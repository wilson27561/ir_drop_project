VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO A2O1A1Ixp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1Ixp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.684 0.272 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.396 0.808 0.468 ;
        RECT 0.216 0.252 0.436 0.324 ;
        RECT 0.216 0.252 0.288 0.468 ;
      LAYER V0 ;
        RECT 0.716 0.396 0.788 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.54 0.98 0.612 ;
        RECT 0.908 0.252 0.98 0.612 ;
        RECT 0.76 0.252 0.98 0.324 ;
      LAYER V0 ;
        RECT 0.908 0.396 0.98 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.54 1.3 0.612 ;
        RECT 1.228 0.316 1.3 0.612 ;
        RECT 1.08 0.396 1.3 0.468 ;
      LAYER V0 ;
        RECT 1.156 0.396 1.228 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 1.444 0.756 ;
        RECT 1.372 0.108 1.444 0.756 ;
        RECT 1.24 0.108 1.444 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.108 1.116 0.18 ;
      RECT 0.396 0.684 0.9 0.756 ;
  END
END A2O1A1Ixp33_ASAP7_6t_fix

MACRO A2O1A1O1Ixp25_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1O1Ixp25_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.412 0.576 0.484 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.272 0.612 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.54 0.872 0.612 ;
        RECT 0.72 0.252 0.872 0.324 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.072 0.54 1.224 0.612 ;
        RECT 1.152 0.108 1.224 0.612 ;
        RECT 1.072 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.504 0.54 1.656 0.612 ;
        RECT 1.584 0.252 1.656 0.612 ;
        RECT 1.504 0.252 1.656 0.324 ;
      LAYER V0 ;
        RECT 1.584 0.4 1.656 0.472 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.476 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.476 0.108 1.548 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.684 1.548 0.756 ;
      RECT 0.396 0.108 0.9 0.18 ;
      RECT 0.18 0.684 0.684 0.756 ;
  END
END A2O1A1O1Ixp25_ASAP7_6t_fix

MACRO AND2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.584 ;
        RECT 0.288 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.392 0.576 0.464 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.36 0.612 ;
        RECT 0.288 0.424 0.36 0.612 ;
        RECT 0.072 0.284 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.288 0.468 0.36 0.54 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.828 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.288 0.684 0.72 0.756 ;
      RECT 0.648 0.108 0.72 0.756 ;
      RECT 0.648 0.396 0.812 0.468 ;
      RECT 0.18 0.108 0.72 0.18 ;
  END
END AND2x1_ASAP7_6t_fix

MACRO AND2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.376 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.24 0.756 ;
        RECT 0.072 0.252 0.224 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 1.08 0.756 ;
        RECT 1.008 0.108 1.08 0.756 ;
        RECT 0.828 0.108 1.08 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 0.72 0.756 ;
      RECT 0.648 0.108 0.72 0.756 ;
      RECT 0.648 0.396 0.812 0.468 ;
      RECT 0.16 0.108 0.72 0.18 ;
  END
END AND2x2_ASAP7_6t_fix

MACRO AND2x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x4_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.008 0.488 ;
        RECT 0.072 0.108 1.008 0.18 ;
        RECT 0.072 0.108 0.144 0.584 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.504 0.596 0.576 ;
        RECT 0.216 0.252 0.488 0.324 ;
        RECT 0.064 0.684 0.288 0.756 ;
        RECT 0.216 0.252 0.288 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.504 0.576 0.576 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.24 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.972 0.756 ;
      RECT 0.9 0.588 0.972 0.756 ;
      RECT 0.72 0.252 0.792 0.756 ;
      RECT 0.9 0.588 1.152 0.66 ;
      RECT 1.08 0.396 1.152 0.66 ;
      RECT 1.08 0.396 1.244 0.468 ;
      RECT 0.612 0.252 0.792 0.324 ;
  END
END AND2x4_ASAP7_6t_fix

MACRO AND2x6_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x6_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.008 0.488 ;
        RECT 0.072 0.108 1.008 0.18 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.504 0.596 0.576 ;
        RECT 0.376 0.252 0.448 0.576 ;
        RECT 0.244 0.252 0.448 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.504 0.576 0.576 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 2.216 0.756 ;
        RECT 1.24 0.108 2.216 0.18 ;
        RECT 1.8 0.108 1.872 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 0.972 0.756 ;
      RECT 0.9 0.588 0.972 0.756 ;
      RECT 0.72 0.252 0.792 0.756 ;
      RECT 0.9 0.588 1.152 0.66 ;
      RECT 1.08 0.396 1.152 0.66 ;
      RECT 1.08 0.396 1.244 0.468 ;
      RECT 0.612 0.252 0.792 0.324 ;
  END
END AND2x6_ASAP7_6t_fix

MACRO AND3x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.364 0.612 ;
        RECT 0.072 0.252 0.252 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5 0.252 0.572 0.468 ;
        RECT 0.392 0.252 0.572 0.324 ;
        RECT 0.392 0.108 0.464 0.324 ;
        RECT 0.06 0.108 0.464 0.18 ;
      LAYER V0 ;
        RECT 0.5 0.344 0.572 0.416 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.54 0.792 0.612 ;
        RECT 0.72 0.328 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 1.044 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.156 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.864 0.396 1.028 0.468 ;
      RECT 0.612 0.108 0.936 0.18 ;
  END
END AND3x1_ASAP7_6t_fix

MACRO AND3x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.264 0.612 ;
        RECT 0.072 0.252 0.264 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.468 ;
        RECT 0.396 0.252 0.576 0.324 ;
        RECT 0.396 0.108 0.468 0.324 ;
        RECT 0.064 0.108 0.468 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.348 0.576 0.42 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.54 0.792 0.612 ;
        RECT 0.72 0.328 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 1.044 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.156 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.864 0.396 1.028 0.468 ;
      RECT 0.612 0.108 0.936 0.18 ;
  END
END AND3x2_ASAP7_6t_fix

MACRO AND3x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x4_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.396 2.776 0.468 ;
        RECT 2.228 0.54 2.52 0.612 ;
        RECT 2.448 0.396 2.52 0.612 ;
      LAYER V0 ;
        RECT 2.556 0.396 2.628 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.396 2.304 0.468 ;
        RECT 1.644 0.54 1.872 0.612 ;
        RECT 1.8 0.396 1.872 0.612 ;
      LAYER V0 ;
        RECT 2.124 0.396 2.196 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.916 0.252 1.764 0.324 ;
        RECT 1.216 0.54 1.52 0.612 ;
        RECT 1.368 0.252 1.44 0.612 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.684 0.92 0.756 ;
        RECT 0.288 0.108 0.92 0.18 ;
        RECT 0.288 0.108 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.684 2.976 0.756 ;
      RECT 2.904 0.108 2.976 0.756 ;
      RECT 1.044 0.396 1.116 0.756 ;
      RECT 0.916 0.396 1.116 0.468 ;
      RECT 2.536 0.108 2.976 0.18 ;
      RECT 1.888 0.252 2.804 0.324 ;
      RECT 1.24 0.108 2.216 0.18 ;
  END
END AND3x4_ASAP7_6t_fix

MACRO AND3x6_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x6_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.236 0.684 3.384 0.756 ;
        RECT 3.312 0.252 3.384 0.756 ;
        RECT 3.236 0.252 3.384 0.324 ;
      LAYER V0 ;
        RECT 3.312 0.396 3.384 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.208 0.54 2.648 0.612 ;
        RECT 2.208 0.396 2.648 0.468 ;
        RECT 2.208 0.396 2.28 0.612 ;
      LAYER V0 ;
        RECT 2.556 0.396 2.628 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.54 1.916 0.612 ;
        RECT 1.584 0.396 1.916 0.468 ;
        RECT 1.584 0.252 1.656 0.612 ;
        RECT 1.256 0.252 1.656 0.324 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 2.976 0.54 3.072 0.912 ;
        RECT 2.544 0.54 2.64 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 1.352 0.18 ;
        RECT 0.072 0.684 1.332 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.44 0.684 2.844 0.756 ;
      RECT 2.772 0.252 2.844 0.756 ;
      RECT 1.44 0.396 1.512 0.756 ;
      RECT 1.152 0.396 1.512 0.468 ;
      RECT 2.772 0.252 3.06 0.324 ;
      RECT 1.908 0.252 2.628 0.324 ;
      RECT 1.908 0.108 1.98 0.324 ;
      RECT 1.584 0.108 1.98 0.18 ;
      RECT 2.34 0.108 3.296 0.18 ;
  END
END AND3x6_ASAP7_6t_fix

MACRO AND4x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.54 0.576 0.612 ;
        RECT 0.504 0.412 0.576 0.612 ;
        RECT 0.288 0.252 0.436 0.324 ;
        RECT 0.288 0.252 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.412 0.576 0.484 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.444 ;
        RECT 0.632 0.252 0.792 0.324 ;
        RECT 0.632 0.108 0.704 0.324 ;
        RECT 0.556 0.108 0.704 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.352 0.792 0.424 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.892 0.256 1.04 0.328 ;
        RECT 0.828 0.54 1.008 0.612 ;
        RECT 0.936 0.256 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.392 1.008 0.464 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3 0.608 1.448 0.756 ;
        RECT 1.3 0.108 1.448 0.256 ;
        RECT 1.368 0.108 1.44 0.756 ;
      LAYER V0 ;
        RECT 1.368 0.536 1.44 0.608 ;
        RECT 1.368 0.256 1.44 0.328 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 1.224 0.756 ;
      RECT 1.152 0.108 1.224 0.756 ;
      RECT 0.828 0.108 1.224 0.18 ;
  END
END AND4x1_ASAP7_6t_fix

MACRO AND4x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.54 1.008 0.612 ;
        RECT 0.936 0.328 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.396 0.576 0.468 ;
        RECT 0.288 0.28 0.36 0.584 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.488 ;
        RECT 0.532 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.24 0.756 ;
        RECT 0.072 0.292 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.512 0.756 ;
        RECT 1.44 0.108 1.512 0.756 ;
        RECT 1.26 0.108 1.512 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 1.152 0.756 ;
      RECT 1.08 0.108 1.152 0.756 ;
      RECT 1.08 0.396 1.224 0.468 ;
      RECT 0.16 0.108 1.152 0.18 ;
  END
END AND4x2_ASAP7_6t_fix

MACRO AND4x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x4_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.224 0.612 ;
        RECT 0.072 0.252 0.224 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.424 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.4 0.576 0.472 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.252 0.796 0.4 ;
        RECT 0.72 0.252 0.792 0.584 ;
      LAYER V0 ;
        RECT 0.72 0.412 0.792 0.484 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.868 0.252 1.016 0.4 ;
        RECT 0.936 0.252 1.008 0.584 ;
      LAYER V0 ;
        RECT 0.936 0.412 1.008 0.484 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.764 0.756 ;
        RECT 1.26 0.108 1.764 0.18 ;
        RECT 1.584 0.108 1.656 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 1.16 0.756 ;
      RECT 1.088 0.108 1.16 0.756 ;
      RECT 1.088 0.396 1.26 0.468 ;
      RECT 0.18 0.108 1.16 0.18 ;
  END
END AND4x4_ASAP7_6t_fix

MACRO AND4x6_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4x6_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.224 0.612 ;
        RECT 0.072 0.252 0.224 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.424 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.4 0.576 0.472 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.252 0.796 0.4 ;
        RECT 0.72 0.252 0.792 0.584 ;
      LAYER V0 ;
        RECT 0.72 0.412 0.792 0.484 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.868 0.252 1.016 0.4 ;
        RECT 0.936 0.252 1.008 0.584 ;
      LAYER V0 ;
        RECT 0.936 0.412 1.008 0.484 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 2.196 0.756 ;
        RECT 1.26 0.108 2.196 0.18 ;
        RECT 1.8 0.108 1.872 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 1.16 0.756 ;
      RECT 1.088 0.108 1.16 0.756 ;
      RECT 1.088 0.396 1.26 0.468 ;
      RECT 0.18 0.108 1.16 0.18 ;
  END
END AND4x6_ASAP7_6t_fix

MACRO AND5x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.224 0.612 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.108 0.576 0.448 ;
        RECT 0.424 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.356 0.576 0.428 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.64 0.54 0.792 0.612 ;
        RECT 0.72 0.416 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.44 0.792 0.512 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.448 ;
        RECT 0.852 0.252 1.008 0.324 ;
      LAYER V0 ;
        RECT 0.936 0.356 1.008 0.428 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.068 0.54 1.224 0.612 ;
        RECT 1.152 0.328 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.236 1.656 0.628 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.684 1.44 0.756 ;
      RECT 1.368 0.108 1.44 0.756 ;
      RECT 1.044 0.108 1.44 0.18 ;
  END
END AND5x1_ASAP7_6t_fix

MACRO AND5x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.36 0.18 ;
        RECT 0.072 0.54 0.224 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.424 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.444 0.576 0.516 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.44 ;
        RECT 0.64 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.368 0.792 0.44 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.732 0.54 1.008 0.612 ;
        RECT 0.936 0.424 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.444 1.008 0.516 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.532 ;
        RECT 0.928 0.252 1.224 0.324 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.684 1.728 0.756 ;
        RECT 1.656 0.108 1.728 0.756 ;
        RECT 1.476 0.108 1.728 0.18 ;
      LAYER V0 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.684 1.368 0.756 ;
      RECT 1.296 0.108 1.368 0.756 ;
      RECT 1.296 0.396 1.46 0.468 ;
      RECT 1.044 0.108 1.368 0.18 ;
  END
END AND5x2_ASAP7_6t_fix

MACRO AO211x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211x2_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.368 0.612 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.496 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.496 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.4 0.792 0.472 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.656 0.468 ;
        RECT 0.936 0.252 1.096 0.608 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 0.252 2.592 0.492 ;
        RECT 1.976 0.252 2.592 0.324 ;
      LAYER V0 ;
        RECT 2.52 0.396 2.592 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 0.816 -0.048 1.128 0.216 ;
        RECT 0.816 -0.048 1.012 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.684 3.384 0.756 ;
        RECT 3.312 0.108 3.384 0.756 ;
        RECT 2.968 0.108 3.384 0.18 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.104 0.684 2.736 0.756 ;
      RECT 2.664 0.108 2.736 0.756 ;
      RECT 2.664 0.396 2.972 0.468 ;
      RECT 0.396 0.108 2.736 0.18 ;
      RECT 1.24 0.54 2.412 0.612 ;
      RECT 0.18 0.684 1.572 0.756 ;
  END
END AO211x2_ASAP7_6t_fix

MACRO AO21x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.22 0.256 ;
        RECT 0.064 0.54 0.212 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 0.568 0.468 ;
        RECT 0.32 0.108 0.488 0.18 ;
        RECT 0.36 0.108 0.432 0.468 ;
      LAYER V0 ;
        RECT 0.496 0.396 0.568 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.692 0.396 0.912 0.468 ;
        RECT 0.84 0.252 0.912 0.468 ;
        RECT 0.692 0.252 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.748 0.396 0.82 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.928 0.684 1.224 0.756 ;
        RECT 1.152 0.136 1.224 0.756 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.336 0.54 1.068 0.612 ;
      RECT 0.996 0.108 1.068 0.612 ;
      RECT 0.612 0.108 1.068 0.18 ;
      RECT 0.18 0.684 0.704 0.756 ;
  END
END AO21x1_ASAP7_6t_fix

MACRO AO21x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.252 0.612 ;
        RECT 0.072 0.136 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 0.576 0.468 ;
        RECT 0.36 0.108 0.432 0.468 ;
        RECT 0.252 0.108 0.432 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.7 0.396 0.888 0.468 ;
        RECT 0.816 0.28 0.888 0.468 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.92 0.684 1.296 0.756 ;
        RECT 1.224 0.276 1.296 0.756 ;
        RECT 1.104 0.276 1.296 0.348 ;
        RECT 1.104 0.152 1.176 0.348 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.104 0.18 1.176 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.54 1.032 0.612 ;
      RECT 0.96 0.108 1.032 0.612 ;
      RECT 0.612 0.108 1.032 0.18 ;
      RECT 0.18 0.684 0.704 0.756 ;
  END
END AO21x2_ASAP7_6t_fix

MACRO AO221x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.54 1.228 0.612 ;
        RECT 1.08 0.324 1.152 0.612 ;
        RECT 0.936 0.324 1.152 0.396 ;
      LAYER V0 ;
        RECT 0.936 0.324 1.008 0.396 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.62 0.684 1.768 0.756 ;
        RECT 1.62 0.54 1.692 0.756 ;
        RECT 1.368 0.54 1.692 0.612 ;
        RECT 1.368 0.252 1.528 0.324 ;
        RECT 1.368 0.252 1.44 0.612 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.464 0.216 0.612 ;
        RECT 0.072 0.24 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.392 0.144 0.464 ;
    END
  END B1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.54 0.868 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.504 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.324 0.792 0.396 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.216 ;
        RECT 0.6 -0.048 0.696 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.908 0.684 2.088 0.756 ;
        RECT 2.016 0.108 2.088 0.756 ;
        RECT 1.908 0.108 2.088 0.18 ;
      LAYER V0 ;
        RECT 1.908 0.684 1.98 0.756 ;
        RECT 1.908 0.108 1.98 0.18 ;
    END
  END Y
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.308 0.396 0.648 0.468 ;
      LAYER M1 ;
        RECT 0.46 0.396 0.62 0.468 ;
      LAYER V1 ;
        RECT 0.504 0.396 0.576 0.468 ;
      LAYER V0 ;
        RECT 0.528 0.396 0.6 0.468 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 0.288 0.54 0.508 0.612 ;
      RECT 0.288 0.108 0.36 0.612 ;
      RECT 1.736 0.108 1.808 0.46 ;
      RECT 0.288 0.108 1.808 0.18 ;
      RECT 0.828 0.684 1.496 0.756 ;
      RECT 0.072 0.684 0.684 0.756 ;
  END
END AO221x1_ASAP7_6t_fix

MACRO AO221x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.54 1.228 0.612 ;
        RECT 1.08 0.324 1.152 0.612 ;
        RECT 0.936 0.324 1.152 0.396 ;
      LAYER V0 ;
        RECT 0.936 0.324 1.008 0.396 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.62 0.684 1.768 0.756 ;
        RECT 1.62 0.54 1.692 0.756 ;
        RECT 1.368 0.54 1.692 0.612 ;
        RECT 1.368 0.252 1.528 0.324 ;
        RECT 1.368 0.252 1.44 0.612 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.464 0.216 0.612 ;
        RECT 0.072 0.24 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.392 0.144 0.464 ;
    END
  END B1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.54 0.868 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.504 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.324 0.792 0.396 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.216 ;
        RECT 0.6 -0.048 0.696 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.908 0.684 2.304 0.756 ;
        RECT 2.232 0.108 2.304 0.756 ;
        RECT 1.908 0.108 2.304 0.18 ;
      LAYER V0 ;
        RECT 1.908 0.684 1.98 0.756 ;
        RECT 1.908 0.108 1.98 0.18 ;
    END
  END Y
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.308 0.396 0.648 0.468 ;
      LAYER M1 ;
        RECT 0.46 0.396 0.62 0.468 ;
      LAYER V1 ;
        RECT 0.504 0.396 0.576 0.468 ;
      LAYER V0 ;
        RECT 0.528 0.396 0.6 0.468 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 0.288 0.54 0.508 0.612 ;
      RECT 0.288 0.108 0.36 0.612 ;
      RECT 1.736 0.108 1.808 0.46 ;
      RECT 0.288 0.108 1.808 0.18 ;
      RECT 0.828 0.684 1.496 0.756 ;
      RECT 0.072 0.684 0.684 0.756 ;
  END
END AO221x2_ASAP7_6t_fix

MACRO AO222x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.776 0.396 2.088 0.468 ;
        RECT 1.776 0.252 2.084 0.324 ;
        RECT 1.776 0.252 1.848 0.468 ;
      LAYER V0 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.54 2.544 0.612 ;
        RECT 2.232 0.28 2.304 0.612 ;
      LAYER V0 ;
        RECT 2.232 0.388 2.304 0.46 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.676 0.468 ;
        RECT 1.368 0.252 1.676 0.324 ;
        RECT 1.368 0.252 1.44 0.468 ;
      LAYER V0 ;
        RECT 1.44 0.396 1.512 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.252 1.236 0.324 ;
        RECT 1.004 0.54 1.152 0.612 ;
        RECT 1.08 0.252 1.152 0.612 ;
      LAYER V0 ;
        RECT 1.08 0.388 1.152 0.46 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.272 0.612 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 0.732 0.468 ;
        RECT 0.504 0.252 0.576 0.468 ;
        RECT 0.424 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.576 0.396 0.648 0.468 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 0.684 2.736 0.756 ;
        RECT 2.664 0.188 2.736 0.756 ;
      LAYER V0 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.664 0.188 2.736 0.26 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.54 0.904 0.612 ;
      RECT 0.832 0.108 0.904 0.612 ;
      RECT 2.388 0.388 2.556 0.46 ;
      RECT 2.388 0.108 2.46 0.46 ;
      RECT 0.396 0.108 2.46 0.18 ;
      RECT 1.8 0.684 2.196 0.756 ;
      RECT 1.8 0.54 1.872 0.756 ;
      RECT 1.28 0.54 1.872 0.612 ;
      RECT 0.18 0.684 1.548 0.756 ;
  END
END AO222x1_ASAP7_6t_fix

MACRO AO222x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.252 1.948 0.324 ;
        RECT 1.8 0.252 1.872 0.492 ;
      LAYER V0 ;
        RECT 1.8 0.4 1.872 0.472 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.54 2.312 0.612 ;
        RECT 2.016 0.38 2.088 0.612 ;
      LAYER V0 ;
        RECT 2.016 0.4 2.088 0.472 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.416 0.252 1.7 0.324 ;
        RECT 1.324 0.396 1.488 0.468 ;
        RECT 1.416 0.252 1.488 0.468 ;
      LAYER V0 ;
        RECT 1.344 0.396 1.416 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.932 0.252 1.232 0.324 ;
        RECT 0.932 0.252 1.08 0.38 ;
        RECT 0.932 0.252 1.004 0.472 ;
      LAYER V0 ;
        RECT 0.932 0.38 1.004 0.452 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.476 ;
        RECT 0.496 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.38 0.792 0.452 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 2.544 0.54 2.64 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 2.544 -0.048 2.64 0.324 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.228 0.684 2.736 0.756 ;
        RECT 2.664 0.108 2.736 0.756 ;
        RECT 2.34 0.108 2.736 0.18 ;
        RECT 2.34 0.108 2.412 0.272 ;
      LAYER V0 ;
        RECT 2.34 0.684 2.412 0.756 ;
        RECT 2.34 0.18 2.412 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.324 0.54 0.648 0.612 ;
      RECT 0.324 0.108 0.396 0.612 ;
      RECT 2.196 0.396 2.412 0.468 ;
      RECT 2.196 0.108 2.268 0.468 ;
      RECT 0.324 0.108 2.268 0.18 ;
      RECT 1.584 0.684 2.088 0.756 ;
      RECT 1.584 0.54 1.656 0.756 ;
      RECT 1.048 0.54 1.656 0.612 ;
      RECT 0.376 0.684 1.352 0.756 ;
  END
END AO222x2_ASAP7_6t_fix

MACRO AO22x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.488 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 0.596 0.468 ;
        RECT 0.284 0.54 0.432 0.612 ;
        RECT 0.36 0.252 0.432 0.612 ;
        RECT 0.284 0.252 0.432 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.684 1.452 0.756 ;
        RECT 1.296 0.324 1.368 0.756 ;
        RECT 0.936 0.324 1.368 0.396 ;
      LAYER V0 ;
        RECT 0.936 0.324 1.008 0.396 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.44 ;
        RECT 0.572 0.252 0.792 0.324 ;
        RECT 0.572 0.108 0.644 0.324 ;
        RECT 0.38 0.108 0.644 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.332 0.792 0.404 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.672 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.44 0.108 1.512 0.468 ;
      RECT 0.828 0.108 1.512 0.18 ;
      RECT 0.18 0.684 1.116 0.756 ;
  END
END AO22x1_ASAP7_6t_fix

MACRO AO22x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.404 0.18 ;
        RECT 0.072 0.396 0.296 0.468 ;
        RECT 0.072 0.54 0.292 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.224 0.396 0.296 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.252 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.384 0.576 0.456 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.448 0.756 ;
        RECT 1.22 0.396 1.44 0.468 ;
        RECT 1.368 0.252 1.44 0.468 ;
        RECT 1.144 0.252 1.44 0.324 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.252 1.332 0.324 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.084 0.468 ;
        RECT 0.936 0.252 1.008 0.468 ;
        RECT 0.696 0.252 1.008 0.324 ;
        RECT 0.696 0.252 0.768 0.476 ;
      LAYER V0 ;
        RECT 0.696 0.384 0.768 0.456 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.684 2.088 0.756 ;
        RECT 2.016 0.108 2.088 0.756 ;
        RECT 1.692 0.108 2.088 0.18 ;
      LAYER V0 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.832 0.54 1.584 0.612 ;
      RECT 1.512 0.108 1.584 0.612 ;
      RECT 1.512 0.396 1.676 0.468 ;
      RECT 0.544 0.108 1.584 0.18 ;
      RECT 0.18 0.684 1.136 0.756 ;
  END
END AO22x2_ASAP7_6t_fix

MACRO AO31x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31x1_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 0.54 2.672 0.612 ;
        RECT 2.52 0.252 2.672 0.324 ;
        RECT 2.52 0.252 2.592 0.612 ;
        RECT 2.024 0.396 2.592 0.468 ;
      LAYER V0 ;
        RECT 2.128 0.396 2.2 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3 0.396 1.9 0.468 ;
        RECT 1.3 0.252 1.372 0.468 ;
        RECT 1.224 0.252 1.372 0.324 ;
      LAYER V0 ;
        RECT 1.692 0.396 1.764 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.22 0.612 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.576 0.396 0.9 0.468 ;
        RECT 0.428 0.54 0.648 0.612 ;
        RECT 0.576 0.252 0.648 0.612 ;
        RECT 0.428 0.252 0.648 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.396 0.9 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.988 0.684 3.168 0.756 ;
        RECT 3.096 0.108 3.168 0.756 ;
        RECT 2.988 0.108 3.168 0.18 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.32 0.684 2.888 0.756 ;
      RECT 2.816 0.108 2.888 0.756 ;
      RECT 2.32 0.54 2.392 0.756 ;
      RECT 0.828 0.54 2.392 0.612 ;
      RECT 1.044 0.252 1.116 0.612 ;
      RECT 2.816 0.396 2.996 0.468 ;
      RECT 0.808 0.252 1.116 0.324 ;
      RECT 2.124 0.108 2.888 0.18 ;
      RECT 1.496 0.252 2.396 0.324 ;
      RECT 0.16 0.684 2.196 0.756 ;
      RECT 0.396 0.108 1.764 0.18 ;
  END
END AO31x1_ASAP7_6t_fix

MACRO AO31x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31x2_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 0.54 2.672 0.612 ;
        RECT 2.52 0.252 2.672 0.324 ;
        RECT 2.52 0.252 2.592 0.612 ;
        RECT 2.024 0.396 2.592 0.468 ;
      LAYER V0 ;
        RECT 2.128 0.396 2.2 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.3 0.396 1.9 0.468 ;
        RECT 1.3 0.252 1.372 0.468 ;
        RECT 1.224 0.252 1.372 0.324 ;
      LAYER V0 ;
        RECT 1.692 0.396 1.764 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.22 0.612 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.576 0.396 0.9 0.468 ;
        RECT 0.428 0.54 0.648 0.612 ;
        RECT 0.576 0.252 0.648 0.612 ;
        RECT 0.428 0.252 0.648 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.396 0.9 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.988 0.684 3.384 0.756 ;
        RECT 3.312 0.108 3.384 0.756 ;
        RECT 2.988 0.108 3.384 0.18 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.32 0.684 2.888 0.756 ;
      RECT 2.816 0.108 2.888 0.756 ;
      RECT 2.32 0.54 2.392 0.756 ;
      RECT 0.828 0.54 2.392 0.612 ;
      RECT 1.044 0.252 1.116 0.612 ;
      RECT 2.816 0.396 2.996 0.468 ;
      RECT 0.828 0.252 1.116 0.324 ;
      RECT 2.124 0.108 2.888 0.18 ;
      RECT 1.496 0.252 2.396 0.324 ;
      RECT 0.16 0.684 2.196 0.756 ;
      RECT 0.396 0.108 1.764 0.18 ;
  END
END AO31x2_ASAP7_6t_fix

MACRO AO322x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO322x2_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.42 0.54 0.568 0.612 ;
        RECT 0.496 0.252 0.568 0.612 ;
        RECT 0.42 0.252 0.568 0.324 ;
      LAYER V0 ;
        RECT 0.496 0.34 0.568 0.412 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.532 0.468 ;
        RECT 1.34 0.108 1.508 0.18 ;
        RECT 1.368 0.108 1.44 0.468 ;
      LAYER V0 ;
        RECT 1.368 0.292 1.44 0.364 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.048 0.252 1.196 0.324 ;
        RECT 0.956 0.38 1.12 0.452 ;
        RECT 1.048 0.252 1.12 0.452 ;
      LAYER V0 ;
        RECT 0.976 0.38 1.048 0.452 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.108 1.872 0.44 ;
        RECT 1.632 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.8 0.328 1.872 0.4 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.108 2.432 0.18 ;
        RECT 2.016 0.108 2.088 0.44 ;
      LAYER V0 ;
        RECT 2.016 0.328 2.088 0.4 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.536 0.684 3.168 0.756 ;
        RECT 3.096 0.108 3.168 0.756 ;
        RECT 2.556 0.108 3.168 0.18 ;
      LAYER V0 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Y
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.5 0.396 0.832 0.468 ;
      LAYER M1 ;
        RECT 0.684 0.396 0.832 0.468 ;
      LAYER V1 ;
        RECT 0.728 0.396 0.8 0.468 ;
      LAYER V0 ;
        RECT 0.716 0.396 0.788 0.468 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 1.656 0.54 2.44 0.612 ;
      RECT 2.368 0.392 2.44 0.612 ;
      RECT 2.368 0.392 2.736 0.464 ;
      RECT 0.376 0.684 0.9 0.756 ;
      RECT 0.68 0.54 0.752 0.756 ;
      RECT 0.68 0.54 1.308 0.612 ;
      RECT 1.024 0.684 2 0.756 ;
      RECT 0.504 0.108 1.116 0.18 ;
  END
END AO322x2_ASAP7_6t_fix

MACRO AO32x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.864 0.108 1.136 0.18 ;
        RECT 0.864 0.396 1.012 0.468 ;
        RECT 0.864 0.108 0.936 0.468 ;
      LAYER V0 ;
        RECT 0.94 0.396 1.012 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.54 1.052 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.392 0.792 0.464 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.384 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.396 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.412 0.576 0.484 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.136 0.396 1.508 0.468 ;
        RECT 1.436 0.252 1.508 0.468 ;
        RECT 1.288 0.252 1.508 0.324 ;
      LAYER V0 ;
        RECT 1.156 0.396 1.228 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.684 1.872 0.756 ;
        RECT 1.8 0.136 1.872 0.756 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.264 0.756 ;
        RECT 0.072 0.248 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.544 0.144 0.616 ;
        RECT 0.072 0.248 0.144 0.32 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.288 0.54 1.652 0.612 ;
      RECT 1.58 0.108 1.652 0.612 ;
      RECT 1.26 0.108 1.652 0.18 ;
      RECT 0.22 0.108 0.292 0.464 ;
      RECT 0.22 0.108 0.684 0.18 ;
      RECT 0.512 0.684 1.568 0.756 ;
  END
END AO32x1_ASAP7_6t_fix

MACRO AO32x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.224 0.488 ;
        RECT 1.076 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.084 0.612 ;
        RECT 0.936 0.252 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.392 1.008 0.464 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.54 0.792 0.612 ;
        RECT 0.72 0.316 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.412 0.792 0.484 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.136 1.44 0.484 ;
      LAYER V0 ;
        RECT 1.368 0.392 1.44 0.464 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.136 1.872 0.56 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.216 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.468 0.756 ;
        RECT 0.072 0.108 0.468 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.524 0.54 1.688 0.612 ;
      RECT 1.616 0.252 1.688 0.612 ;
      RECT 1.524 0.252 1.688 0.324 ;
      RECT 1.524 0.156 1.596 0.324 ;
      RECT 0.288 0.256 0.36 0.464 ;
      RECT 0.288 0.256 0.648 0.328 ;
      RECT 0.576 0.108 0.648 0.328 ;
      RECT 0.576 0.108 0.9 0.18 ;
      RECT 0.728 0.684 1.784 0.756 ;
  END
END AO32x2_ASAP7_6t_fix

MACRO AO331x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.912 0.108 1.06 0.18 ;
        RECT 0.912 0.108 0.984 0.572 ;
      LAYER V0 ;
        RECT 0.912 0.396 0.984 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.692 0.464 0.84 0.612 ;
        RECT 0.708 0.28 0.78 0.612 ;
      LAYER V0 ;
        RECT 0.708 0.392 0.78 0.464 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.056 0.396 1.22 0.468 ;
        RECT 1.056 0.316 1.128 0.468 ;
      LAYER V0 ;
        RECT 1.128 0.396 1.2 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.32 0.384 1.484 0.456 ;
        RECT 1.32 0.108 1.392 0.456 ;
        RECT 1.244 0.108 1.392 0.18 ;
      LAYER V0 ;
        RECT 1.392 0.384 1.464 0.456 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.608 0.396 1.8 0.468 ;
        RECT 1.728 0.28 1.8 0.468 ;
      LAYER V0 ;
        RECT 1.608 0.396 1.68 0.468 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.872 0.684 2.02 0.756 ;
        RECT 1.872 0.384 1.944 0.756 ;
      LAYER V0 ;
        RECT 1.872 0.404 1.944 0.476 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.272 0.756 ;
        RECT 0.072 0.18 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.492 0.108 1.564 0.252 ;
      RECT 1.492 0.108 1.98 0.18 ;
      RECT 1.692 0.54 1.764 0.684 ;
      RECT 1.22 0.54 1.764 0.612 ;
      RECT 0.22 0.108 0.292 0.468 ;
      RECT 0.22 0.108 0.684 0.18 ;
      RECT 0.456 0.684 1.548 0.756 ;
  END
END AO331x1_ASAP7_6t_fix

MACRO AO331x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.128 0.108 1.2 0.468 ;
        RECT 1.052 0.108 1.2 0.18 ;
      LAYER V0 ;
        RECT 1.128 0.396 1.2 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.924 0.54 1.072 0.612 ;
        RECT 0.924 0.252 0.996 0.612 ;
        RECT 0.712 0.252 0.996 0.324 ;
      LAYER V0 ;
        RECT 0.924 0.396 0.996 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.576 0.54 0.796 0.612 ;
        RECT 0.576 0.396 0.796 0.468 ;
        RECT 0.576 0.396 0.648 0.612 ;
      LAYER V0 ;
        RECT 0.724 0.396 0.796 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.272 0.396 1.436 0.468 ;
        RECT 1.272 0.172 1.344 0.468 ;
      LAYER V0 ;
        RECT 1.344 0.396 1.416 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.536 0.384 1.7 0.456 ;
        RECT 1.536 0.108 1.608 0.456 ;
        RECT 1.46 0.108 1.608 0.18 ;
      LAYER V0 ;
        RECT 1.608 0.384 1.68 0.456 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.824 0.396 1.972 0.468 ;
        RECT 1.9 0.28 1.972 0.468 ;
      LAYER V0 ;
        RECT 1.824 0.396 1.896 0.468 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.084 0.684 2.304 0.756 ;
        RECT 2.084 0.408 2.156 0.756 ;
      LAYER V0 ;
        RECT 2.084 0.408 2.156 0.48 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.684 0.488 0.756 ;
        RECT 0.288 0.252 0.468 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.252 0.468 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.692 0.108 1.764 0.256 ;
      RECT 1.692 0.108 2.196 0.18 ;
      RECT 1.908 0.54 1.98 0.684 ;
      RECT 1.436 0.54 1.98 0.612 ;
      RECT 0.072 0.108 0.144 0.468 ;
      RECT 0.072 0.108 0.9 0.18 ;
      RECT 0.672 0.684 1.764 0.756 ;
  END
END AO331x2_ASAP7_6t_fix

MACRO AO332x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.108 0.98 0.476 ;
        RECT 0.832 0.108 0.98 0.18 ;
      LAYER V0 ;
        RECT 0.908 0.384 0.98 0.456 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.496 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.352 0.792 0.424 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.404 0.396 0.576 0.468 ;
        RECT 0.328 0.684 0.476 0.756 ;
        RECT 0.404 0.396 0.476 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.052 0.396 1.228 0.468 ;
        RECT 1.052 0.136 1.124 0.468 ;
      LAYER V0 ;
        RECT 1.124 0.396 1.196 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.256 1.44 0.44 ;
        RECT 1.296 0.108 1.376 0.328 ;
        RECT 1.228 0.108 1.376 0.18 ;
      LAYER V0 ;
        RECT 1.368 0.348 1.44 0.42 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.136 2.304 0.568 ;
      LAYER V0 ;
        RECT 2.232 0.396 2.304 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.78 0.252 1.988 0.324 ;
        RECT 1.78 0.252 1.852 0.476 ;
      LAYER V0 ;
        RECT 1.78 0.384 1.852 0.456 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.608 0.228 0.756 ;
        RECT 0.072 0.136 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.156 0.144 0.228 ;
    END
  END Y
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.344 0.396 1.692 0.468 ;
      LAYER M1 ;
        RECT 1.6 0.364 1.672 0.476 ;
      LAYER V1 ;
        RECT 1.6 0.396 1.672 0.468 ;
      LAYER V0 ;
        RECT 1.6 0.384 1.672 0.456 ;
    END
  END B3
  OBS
    LAYER M1 ;
      RECT 1.924 0.54 2.16 0.612 ;
      RECT 2.088 0.108 2.16 0.612 ;
      RECT 1.476 0.108 2.16 0.18 ;
      RECT 0.584 0.684 1.116 0.756 ;
      RECT 1.044 0.54 1.116 0.756 ;
      RECT 1.044 0.54 1.548 0.612 ;
      RECT 0.232 0.108 0.304 0.472 ;
      RECT 0.232 0.108 0.684 0.18 ;
      RECT 1.26 0.684 2.224 0.756 ;
  END
END AO332x1_ASAP7_6t_fix

MACRO AO332x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.124 0.108 1.196 0.476 ;
        RECT 1.048 0.108 1.196 0.18 ;
      LAYER V0 ;
        RECT 1.124 0.384 1.196 0.456 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.54 1.008 0.612 ;
        RECT 0.936 0.296 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.352 1.008 0.424 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.468 ;
        RECT 0.62 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.268 0.396 1.444 0.468 ;
        RECT 1.268 0.108 1.416 0.18 ;
        RECT 1.268 0.108 1.34 0.468 ;
      LAYER V0 ;
        RECT 1.34 0.396 1.412 0.468 ;
    END
  END B1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.996 0.252 2.348 0.324 ;
        RECT 1.996 0.252 2.068 0.476 ;
      LAYER V0 ;
        RECT 1.996 0.384 2.068 0.456 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.208 0.684 0.488 0.756 ;
        RECT 0.288 0.252 0.488 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.252 0.468 0.324 ;
    END
  END Y
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.504 0.252 1.74 0.324 ;
      LAYER M1 ;
        RECT 1.564 0.252 1.728 0.324 ;
        RECT 1.584 0.252 1.656 0.44 ;
      LAYER V1 ;
        RECT 1.648 0.252 1.72 0.324 ;
      LAYER V0 ;
        RECT 1.584 0.348 1.656 0.42 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.56 0.396 1.908 0.468 ;
      LAYER M1 ;
        RECT 1.816 0.364 1.888 0.476 ;
      LAYER V1 ;
        RECT 1.816 0.396 1.888 0.468 ;
      LAYER V0 ;
        RECT 1.816 0.384 1.888 0.456 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.14 0.396 2.524 0.468 ;
      LAYER M1 ;
        RECT 2.2 0.396 2.348 0.468 ;
      LAYER V1 ;
        RECT 2.256 0.396 2.328 0.468 ;
      LAYER V0 ;
        RECT 2.276 0.396 2.348 0.468 ;
    END
  END C1
  OBS
    LAYER M1 ;
      RECT 2.12 0.54 2.52 0.612 ;
      RECT 2.448 0.108 2.52 0.612 ;
      RECT 1.692 0.108 2.52 0.18 ;
      RECT 0.8 0.684 1.332 0.756 ;
      RECT 1.26 0.54 1.332 0.756 ;
      RECT 1.26 0.54 1.764 0.612 ;
      RECT 0.072 0.108 0.144 0.468 ;
      RECT 0.072 0.108 0.9 0.18 ;
      RECT 1.476 0.684 2.44 0.756 ;
  END
END AO332x2_ASAP7_6t_fix

MACRO AO333x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.868 0.324 ;
        RECT 0.644 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.4 0.792 0.472 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.492 0.252 0.564 0.492 ;
        RECT 0.416 0.252 0.564 0.324 ;
      LAYER V0 ;
        RECT 0.492 0.4 0.564 0.472 ;
    END
  END A3
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.34 0.108 1.412 0.44 ;
        RECT 1.264 0.108 1.412 0.18 ;
      LAYER V0 ;
        RECT 1.34 0.344 1.412 0.416 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.124 0.252 1.196 0.476 ;
        RECT 1.052 0.108 1.124 0.324 ;
        RECT 0.976 0.108 1.124 0.18 ;
      LAYER V0 ;
        RECT 1.124 0.384 1.196 0.456 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.304 0.108 2.524 0.18 ;
        RECT 2.304 0.108 2.376 0.456 ;
      LAYER V0 ;
        RECT 2.304 0.384 2.376 0.456 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.252 0.756 ;
        RECT 0.072 0.36 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.54 1.232 0.612 ;
      LAYER M1 ;
        RECT 0.892 0.54 1.04 0.612 ;
        RECT 0.936 0.392 1.008 0.612 ;
      LAYER V1 ;
        RECT 0.936 0.54 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.392 1.008 0.464 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.204 0.396 1.66 0.468 ;
      LAYER M1 ;
        RECT 1.512 0.396 1.66 0.468 ;
      LAYER V1 ;
        RECT 1.556 0.396 1.628 0.468 ;
      LAYER V0 ;
        RECT 1.556 0.396 1.628 0.468 ;
    END
  END B1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.784 0.252 2.24 0.324 ;
      LAYER M1 ;
        RECT 2.024 0.252 2.204 0.324 ;
        RECT 2.024 0.252 2.096 0.436 ;
      LAYER V1 ;
        RECT 2.112 0.252 2.184 0.324 ;
      LAYER V0 ;
        RECT 2.024 0.344 2.096 0.416 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.784 0.396 2.24 0.468 ;
      LAYER M1 ;
        RECT 1.784 0.396 1.952 0.468 ;
        RECT 1.88 0.284 1.952 0.468 ;
      LAYER V1 ;
        RECT 1.808 0.396 1.88 0.468 ;
      LAYER V0 ;
        RECT 1.808 0.396 1.88 0.468 ;
    END
  END C3
  OBS
    LAYER M1 ;
      RECT 1.692 0.54 1.764 0.684 ;
      RECT 1.26 0.54 2.236 0.612 ;
      RECT 1.484 0.108 1.556 0.256 ;
      RECT 1.484 0.108 2.024 0.18 ;
      RECT 0.22 0.108 0.292 0.488 ;
      RECT 0.22 0.108 0.72 0.18 ;
      RECT 1.908 0.684 2.412 0.756 ;
      RECT 0.592 0.684 1.548 0.756 ;
  END
END AO333x1_ASAP7_6t_fix

MACRO AO333x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.104 0.54 1.252 0.612 ;
        RECT 1.144 0.252 1.216 0.612 ;
        RECT 1.068 0.252 1.216 0.324 ;
      LAYER V0 ;
        RECT 1.144 0.396 1.216 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.54 1.004 0.612 ;
        RECT 0.932 0.388 1.004 0.612 ;
      LAYER V0 ;
        RECT 0.932 0.408 1.004 0.48 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.564 0.252 0.836 0.324 ;
        RECT 0.564 0.396 0.792 0.468 ;
        RECT 0.564 0.252 0.636 0.468 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.784 0.252 2.052 0.324 ;
        RECT 1.8 0.252 1.872 0.476 ;
      LAYER V0 ;
        RECT 1.8 0.384 1.872 0.456 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.612 0.252 1.684 0.472 ;
        RECT 1.46 0.252 1.684 0.324 ;
      LAYER V0 ;
        RECT 1.612 0.344 1.684 0.416 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.108 1.548 0.18 ;
        RECT 1.288 0.396 1.508 0.468 ;
        RECT 1.288 0.108 1.36 0.468 ;
      LAYER V0 ;
        RECT 1.36 0.396 1.432 0.468 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.592 0.396 2.74 0.612 ;
        RECT 2.668 0.108 2.74 0.612 ;
        RECT 2.364 0.108 2.74 0.18 ;
        RECT 2.436 0.396 2.74 0.468 ;
      LAYER V0 ;
        RECT 2.52 0.396 2.592 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.24 0.252 2.568 0.324 ;
        RECT 2.24 0.252 2.312 0.436 ;
      LAYER V0 ;
        RECT 2.24 0.344 2.312 0.416 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.972 0.396 2.14 0.468 ;
      LAYER V0 ;
        RECT 2.024 0.396 2.096 0.468 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.492 0.756 ;
        RECT 0.42 0.252 0.492 0.756 ;
        RECT 0.26 0.252 0.492 0.324 ;
      LAYER V0 ;
        RECT 0.348 0.252 0.42 0.324 ;
        RECT 0.42 0.54 0.492 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.928 0.54 2 0.684 ;
      RECT 1.928 0.54 2.4 0.612 ;
      RECT 0.088 0.108 0.16 0.488 ;
      RECT 0.088 0.108 0.9 0.18 ;
      RECT 2.124 0.684 2.628 0.756 ;
      RECT 1.672 0.108 2.24 0.18 ;
      RECT 0.808 0.684 1.764 0.756 ;
      RECT 1.42 0.54 1.568 0.612 ;
    LAYER M2 ;
      RECT 1.468 0.54 2.028 0.612 ;
    LAYER V1 ;
      RECT 1.936 0.54 2.008 0.612 ;
      RECT 1.488 0.54 1.56 0.612 ;
  END
END AO333x2_ASAP7_6t_fix

MACRO AO33x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.112 1.008 0.468 ;
        RECT 0.86 0.112 1.008 0.184 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.54 0.868 0.612 ;
        RECT 0.72 0.28 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.384 0.54 0.576 0.612 ;
        RECT 0.504 0.28 0.576 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.388 0.576 0.46 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.54 1.224 0.612 ;
        RECT 1.152 0.396 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.28 0.252 1.532 0.324 ;
        RECT 1.368 0.252 1.44 0.412 ;
      LAYER V0 ;
        RECT 1.368 0.34 1.44 0.412 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.58 0.396 1.728 0.468 ;
        RECT 1.656 0.28 1.728 0.468 ;
      LAYER V0 ;
        RECT 1.58 0.396 1.652 0.468 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.144 0.684 0.488 0.756 ;
        RECT 0.144 0.108 0.216 0.756 ;
        RECT 0.068 0.108 0.216 0.18 ;
      LAYER V0 ;
        RECT 0.144 0.596 0.216 0.668 ;
        RECT 0.144 0.18 0.216 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.692 0.54 1.764 0.684 ;
      RECT 1.324 0.54 1.872 0.612 ;
      RECT 1.8 0.108 1.872 0.612 ;
      RECT 1.476 0.108 1.872 0.18 ;
      RECT 0.288 0.108 0.36 0.452 ;
      RECT 0.288 0.108 0.684 0.18 ;
      RECT 0.612 0.684 1.548 0.756 ;
  END
END AO33x1_ASAP7_6t_fix

MACRO AO33x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8 0.54 1.216 0.612 ;
        RECT 1.144 0.384 1.216 0.612 ;
      LAYER V0 ;
        RECT 1.144 0.384 1.216 0.456 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.888 0.396 1.036 0.468 ;
        RECT 0.888 0.252 0.96 0.468 ;
        RECT 0.648 0.252 0.96 0.324 ;
      LAYER V0 ;
        RECT 0.964 0.396 1.036 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 0.764 0.468 ;
        RECT 0.36 0.54 0.644 0.612 ;
        RECT 0.36 0.396 0.432 0.612 ;
      LAYER V0 ;
        RECT 0.692 0.396 0.764 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.36 0.252 1.432 0.476 ;
        RECT 1.284 0.252 1.432 0.324 ;
      LAYER V0 ;
        RECT 1.36 0.384 1.432 0.456 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.532 0.396 1.732 0.468 ;
        RECT 1.66 0.28 1.732 0.468 ;
      LAYER V0 ;
        RECT 1.588 0.396 1.66 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.948 0.396 2.112 0.468 ;
        RECT 1.948 0.108 2.096 0.18 ;
        RECT 1.948 0.108 2.02 0.468 ;
      LAYER V0 ;
        RECT 2.02 0.396 2.092 0.468 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.684 0.576 0.756 ;
        RECT 0.216 0.252 0.44 0.324 ;
        RECT 0.216 0.252 0.288 0.756 ;
      LAYER V0 ;
        RECT 0.348 0.252 0.42 0.324 ;
        RECT 0.396 0.684 0.468 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.888 0.684 2.108 0.756 ;
      RECT 2.036 0.54 2.108 0.756 ;
      RECT 1.496 0.54 2.108 0.612 ;
      RECT 1.804 0.108 1.876 0.612 ;
      RECT 0.072 0.108 0.144 0.468 ;
      RECT 0.072 0.108 1.876 0.18 ;
      RECT 0.796 0.684 1.764 0.756 ;
  END
END AO33x2_ASAP7_6t_fix

MACRO AOI211x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.976 0.324 ;
        RECT 0.496 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.872 0.468 ;
        RECT 1.8 0.28 1.872 0.468 ;
        RECT 1.368 0.252 1.44 0.468 ;
        RECT 1.144 0.252 1.44 0.324 ;
      LAYER V0 ;
        RECT 1.532 0.396 1.604 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.396 2.304 0.468 ;
        RECT 2.232 0.252 2.304 0.468 ;
        RECT 2.016 0.252 2.304 0.324 ;
      LAYER V0 ;
        RECT 2.124 0.396 2.196 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.076 0.54 2.52 0.612 ;
        RECT 2.448 0.108 2.52 0.612 ;
        RECT 0.364 0.108 2.52 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 1.908 0.108 1.98 0.18 ;
        RECT 2.124 0.54 2.196 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.684 1.224 0.756 ;
      RECT 1.152 0.54 1.224 0.756 ;
      RECT 1.152 0.54 1.796 0.612 ;
      RECT 1.444 0.684 2.432 0.756 ;
  END
END AOI211x1_ASAP7_6t_fix

MACRO AOI211xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5 0.252 1.268 0.324 ;
        RECT 0.504 0.252 0.576 0.408 ;
      LAYER V0 ;
        RECT 0.504 0.336 0.576 0.408 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.252 0.612 ;
        RECT 0.18 0.108 0.252 0.612 ;
        RECT 0.072 0.108 0.252 0.18 ;
      LAYER V0 ;
        RECT 0.18 0.396 0.252 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.996 0.684 1.44 0.756 ;
        RECT 0.996 0.396 1.068 0.756 ;
        RECT 0.7 0.396 1.068 0.468 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.168 0.54 1.44 0.612 ;
        RECT 1.368 0.108 1.44 0.612 ;
        RECT 1.024 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.6 -0.048 0.696 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.324 0.108 0.9 0.18 ;
        RECT 0.324 0.54 0.896 0.612 ;
        RECT 0.324 0.108 0.396 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.54 0.468 0.612 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.684 0.684 0.756 ;
  END
END AOI211xp5_ASAP7_6t_fix

MACRO AOI21x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 1.224 0.468 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.252 1.08 0.324 ;
      LAYER V0 ;
        RECT 0.668 0.252 0.74 0.324 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.54 1.44 0.612 ;
        RECT 1.368 0.32 1.44 0.612 ;
        RECT 0.288 0.396 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.288 0.396 0.36 0.468 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 0.072 0.108 1.656 0.18 ;
        RECT 0.072 0.108 0.144 0.676 ;
      LAYER V0 ;
        RECT 0.072 0.604 0.144 0.676 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.476 0.684 1.548 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 1.352 0.756 ;
  END
END AOI21x1_ASAP7_6t_fix

MACRO AOI21xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.54 0.62 0.612 ;
        RECT 0.216 0.288 0.568 0.36 ;
        RECT 0.216 0.252 0.476 0.36 ;
        RECT 0.216 0.252 0.288 0.612 ;
      LAYER V0 ;
        RECT 0.476 0.288 0.548 0.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.684 0.292 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.288 0.144 0.36 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.416 0.684 0.792 0.756 ;
        RECT 0.72 0.3 0.792 0.756 ;
      LAYER V0 ;
        RECT 0.72 0.3 0.792 0.372 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.008 0.728 ;
        RECT 0.612 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 0.936 0.54 1.008 0.612 ;
    END
  END Y
END AOI21xp33_ASAP7_6t_fix

MACRO AOI21xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.244 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.392 0.576 0.464 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.432 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.54 1.012 0.612 ;
        RECT 0.676 0.252 0.824 0.324 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.392 0.792 0.464 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.008 0.428 ;
        RECT 0.568 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 0.936 0.356 1.008 0.428 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 0.684 0.756 ;
  END
END AOI21xp5_ASAP7_6t_fix

MACRO AOI221x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221x1_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.396 0.944 0.468 ;
        RECT 0.72 0.108 0.792 0.468 ;
        RECT 0.564 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.832 0.396 0.904 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.488 0.612 ;
        RECT 0.072 0.108 0.44 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.396 1.368 0.468 ;
        RECT 1.08 0.252 1.316 0.324 ;
        RECT 1.08 0.252 1.152 0.468 ;
      LAYER V0 ;
        RECT 1.256 0.396 1.328 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.252 2.24 0.324 ;
        RECT 1.672 0.396 2.164 0.468 ;
        RECT 2.092 0.252 2.164 0.468 ;
      LAYER V0 ;
        RECT 1.696 0.396 1.768 0.468 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.364 0.396 2.78 0.468 ;
        RECT 2.364 0.252 2.78 0.324 ;
        RECT 2.156 0.54 2.436 0.612 ;
        RECT 2.364 0.252 2.436 0.612 ;
      LAYER V0 ;
        RECT 2.56 0.396 2.632 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 2.544 -0.048 2.64 0.216 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.56 0.54 2.952 0.612 ;
        RECT 2.88 0.108 2.952 0.612 ;
        RECT 1.044 0.108 2.952 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 2.34 0.108 2.412 0.18 ;
        RECT 2.56 0.54 2.632 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.684 0.9 0.756 ;
      RECT 0.828 0.54 0.9 0.756 ;
      RECT 0.828 0.54 2 0.612 ;
      RECT 1.24 0.684 2.864 0.756 ;
  END
END AOI221x1_ASAP7_6t_fix

MACRO AOI221xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.54 1.556 0.612 ;
        RECT 1.152 0.108 1.428 0.18 ;
        RECT 1.152 0.108 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.68 0.54 1.872 0.612 ;
        RECT 1.8 0.108 1.872 0.612 ;
        RECT 1.552 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.172 0.144 0.54 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.484 0.396 0.792 0.468 ;
        RECT 0.556 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.52 0.396 0.592 0.468 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.892 0.252 1.04 0.324 ;
        RECT 0.828 0.684 1.008 0.756 ;
        RECT 0.936 0.252 1.008 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.216 ;
        RECT 0.6 -0.048 0.696 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.9 0.18 ;
        RECT 0.288 0.54 0.436 0.612 ;
        RECT 0.288 0.108 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.364 0.54 0.436 0.612 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.24 0.684 1.764 0.756 ;
      RECT 0.18 0.684 0.684 0.756 ;
  END
END AOI221xp5_ASAP7_6t_fix

MACRO AOI222xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222xp33_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.136 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.388 0.396 0.792 0.468 ;
        RECT 0.72 0.252 0.792 0.468 ;
        RECT 0.572 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.324 0.792 0.396 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.396 1.684 0.468 ;
        RECT 1.536 0.108 1.684 0.468 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.252 1.464 0.324 ;
        RECT 1.392 0.108 1.464 0.324 ;
        RECT 1.244 0.108 1.464 0.18 ;
        RECT 0.76 0.54 0.98 0.612 ;
        RECT 0.908 0.252 0.98 0.612 ;
      LAYER V0 ;
        RECT 0.908 0.328 0.98 0.4 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.108 2.304 0.18 ;
        RECT 1.8 0.396 2.132 0.468 ;
        RECT 1.8 0.108 1.872 0.468 ;
      LAYER V0 ;
        RECT 1.8 0.284 1.872 0.356 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.684 2.304 0.756 ;
        RECT 2.232 0.28 2.304 0.756 ;
      LAYER V0 ;
        RECT 2.232 0.396 2.304 0.468 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 0.816 -0.048 0.912 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.108 1.116 0.18 ;
        RECT 0.216 0.54 0.636 0.612 ;
        RECT 0.216 0.108 0.288 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.564 0.54 0.636 0.612 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.092 0.54 1.98 0.612 ;
      RECT 0.396 0.684 1.352 0.756 ;
  END
END AOI222xp33_ASAP7_6t_fix

MACRO AOI22x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.148 0.252 1.74 0.324 ;
      LAYER V0 ;
        RECT 1.648 0.252 1.72 0.324 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.124 0.396 1.916 0.468 ;
      LAYER V0 ;
        RECT 1.124 0.396 1.196 0.468 ;
        RECT 1.844 0.396 1.916 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.396 0.812 0.468 ;
        RECT 0.612 0.252 0.684 0.468 ;
        RECT 0.2 0.252 0.684 0.324 ;
        RECT 0.2 0.108 0.272 0.324 ;
        RECT 0.064 0.108 0.272 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 1.008 0.612 ;
        RECT 0.936 0.372 1.008 0.612 ;
        RECT 0.072 0.396 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.144 0.54 2.088 0.612 ;
        RECT 2.016 0.108 2.088 0.612 ;
        RECT 0.396 0.108 2.088 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 1.26 0.54 1.332 0.612 ;
        RECT 1.692 0.54 1.764 0.612 ;
        RECT 1.908 0.108 1.98 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 2 0.756 ;
  END
END AOI22x1_ASAP7_6t_fix

MACRO AOI22xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.136 0.144 0.584 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.108 0.576 0.372 ;
        RECT 0.288 0.108 0.576 0.18 ;
        RECT 0.288 0.108 0.36 0.584 ;
      LAYER V0 ;
        RECT 0.504 0.3 0.576 0.372 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.292 0.684 1.44 0.756 ;
        RECT 1.368 0.136 1.44 0.756 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.396 1.084 0.468 ;
        RECT 0.648 0.252 0.868 0.324 ;
        RECT 0.484 0.54 0.72 0.612 ;
        RECT 0.648 0.252 0.72 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.844 0.54 1.256 0.612 ;
        RECT 1.184 0.108 1.256 0.612 ;
        RECT 0.828 0.108 1.256 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 0.864 0.54 0.936 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.064 0.684 1.116 0.756 ;
  END
END AOI22xp33_ASAP7_6t_fix

MACRO AOI22xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.22 0.612 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.392 0.576 0.464 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.136 1.224 0.584 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.392 0.812 0.464 ;
        RECT 0.648 0.108 0.72 0.464 ;
        RECT 0.432 0.108 0.72 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.392 0.792 0.464 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.708 0.54 1.008 0.612 ;
        RECT 0.936 0.108 1.008 0.612 ;
        RECT 0.828 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 0.86 0.54 0.932 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 1.136 0.756 ;
  END
END AOI22xp5_ASAP7_6t_fix

MACRO AOI311xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI311xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.868 0.324 ;
        RECT 0.72 0.252 0.792 0.576 ;
      LAYER V0 ;
        RECT 0.72 0.408 0.792 0.48 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.108 0.576 0.48 ;
        RECT 0.428 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.408 0.576 0.48 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.396 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.084 0.612 ;
        RECT 0.936 0.38 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.408 1.008 0.48 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.224 0.252 1.296 0.56 ;
        RECT 1.148 0.252 1.296 0.324 ;
      LAYER V0 ;
        RECT 1.224 0.408 1.296 0.48 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 0.792 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 0.936 0.756 ;
  END
END AOI311xp33_ASAP7_6t_fix

MACRO AOI31xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.396 0.976 0.468 ;
        RECT 0.72 0.54 0.94 0.612 ;
        RECT 0.72 0.108 0.792 0.612 ;
        RECT 0.424 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.792 0.396 0.864 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.288 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.3 0.18 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.284 0.396 1.484 0.468 ;
        RECT 1.024 0.684 1.356 0.756 ;
        RECT 1.284 0.252 1.356 0.756 ;
        RECT 1.024 0.252 1.356 0.324 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.024 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 1.476 0.684 1.548 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.9 0.756 ;
  END
END AOI31xp33_ASAP7_6t_fix

MACRO AOI31xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31xp67_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.536 0.252 2.736 0.612 ;
        RECT 2.12 0.396 2.736 0.468 ;
      LAYER V0 ;
        RECT 2.12 0.396 2.192 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.28 0.396 1.764 0.468 ;
        RECT 1.28 0.252 1.352 0.468 ;
        RECT 1.204 0.252 1.352 0.324 ;
      LAYER V0 ;
        RECT 1.692 0.396 1.764 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.38 0.612 ;
        RECT 0.072 0.244 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 0.9 0.468 ;
        RECT 0.504 0.252 0.576 0.468 ;
        RECT 0.28 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.396 0.9 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.56 0.828 2.632 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.56 -0.036 2.632 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.34 0.684 2.632 0.756 ;
        RECT 2.34 0.54 2.412 0.756 ;
        RECT 0.828 0.54 2.412 0.612 ;
        RECT 1.008 0.252 1.08 0.612 ;
        RECT 0.828 0.252 1.08 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.54 0.9 0.612 ;
        RECT 0.828 0.252 0.9 0.324 ;
        RECT 2.56 0.684 2.632 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.124 0.108 2.632 0.18 ;
      RECT 1.476 0.252 2.412 0.324 ;
      RECT 0.18 0.684 2.196 0.756 ;
      RECT 0.396 0.108 1.764 0.18 ;
  END
END AOI31xp67_ASAP7_6t_fix

MACRO AOI321xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI321xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.484 ;
        RECT 0.532 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.392 0.792 0.464 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 0.58 0.468 ;
        RECT 0.36 0.108 0.432 0.468 ;
        RECT 0.28 0.108 0.432 0.18 ;
      LAYER V0 ;
        RECT 0.508 0.396 0.58 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.396 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.452 ;
        RECT 1.076 0.252 1.224 0.324 ;
      LAYER V0 ;
        RECT 1.152 0.324 1.224 0.396 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.336 0.396 1.484 0.468 ;
        RECT 1.368 0.28 1.44 0.468 ;
      LAYER V0 ;
        RECT 1.368 0.324 1.44 0.396 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.54 1.084 0.612 ;
        RECT 0.936 0.372 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.392 1.008 0.464 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.54 1.656 0.612 ;
        RECT 1.584 0.108 1.656 0.612 ;
        RECT 0.612 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.26 0.54 1.332 0.612 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.684 1.548 0.756 ;
      RECT 0.396 0.684 0.9 0.756 ;
  END
END AOI321xp33_ASAP7_6t_fix

MACRO AOI322xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI322xp5_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.632 0.396 0.78 0.468 ;
        RECT 0.632 0.108 0.704 0.468 ;
        RECT 0.532 0.108 0.704 0.18 ;
      LAYER V0 ;
        RECT 0.708 0.396 0.78 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.912 0.256 0.984 0.44 ;
        RECT 0.776 0.108 0.944 0.256 ;
        RECT 0.84 0.256 0.984 0.324 ;
      LAYER V0 ;
        RECT 0.912 0.348 0.984 0.42 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.54 1.448 0.612 ;
        RECT 1.296 0.252 1.448 0.324 ;
        RECT 1.296 0.252 1.368 0.612 ;
        RECT 1.088 0.396 1.368 0.468 ;
      LAYER V0 ;
        RECT 1.164 0.396 1.236 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.476 0.32 0.548 0.484 ;
        RECT 0.36 0.32 0.548 0.392 ;
        RECT 0.36 0.108 0.432 0.392 ;
        RECT 0.284 0.108 0.432 0.256 ;
      LAYER V0 ;
        RECT 0.476 0.392 0.548 0.464 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.28 0.612 ;
        RECT 0.064 0.108 0.212 0.256 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.216 2.304 0.54 ;
      LAYER V0 ;
        RECT 2.232 0.396 2.304 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.728 0.252 1.88 0.324 ;
        RECT 1.572 0.54 1.8 0.612 ;
        RECT 1.728 0.252 1.8 0.612 ;
        RECT 1.564 0.396 1.8 0.468 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.936 0.54 2.16 0.612 ;
        RECT 2.088 0.108 2.16 0.612 ;
        RECT 1.044 0.108 2.16 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 1.956 0.54 2.028 0.612 ;
        RECT 2.088 0.18 2.16 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.156 0.684 0.684 0.756 ;
      RECT 0.612 0.54 0.684 0.756 ;
      RECT 0.612 0.54 1.12 0.612 ;
      RECT 0.808 0.684 2.196 0.756 ;
  END
END AOI322xp5_ASAP7_6t_fix

MACRO AOI32x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.54 1.304 0.612 ;
        RECT 1.152 0.34 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.404 1.224 0.476 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.108 1.664 0.18 ;
        RECT 1.368 0.108 1.44 0.436 ;
      LAYER V0 ;
        RECT 1.368 0.344 1.44 0.416 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.684 1.872 0.756 ;
        RECT 1.8 0.252 1.872 0.756 ;
        RECT 1.576 0.252 1.872 0.324 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.452 ;
        RECT 0.368 0.252 1.008 0.324 ;
        RECT 0.268 0.388 0.44 0.46 ;
        RECT 0.368 0.252 0.44 0.46 ;
      LAYER V0 ;
        RECT 0.268 0.388 0.34 0.46 ;
        RECT 0.936 0.38 1.008 0.452 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.152 0.108 1.152 0.18 ;
      LAYER M1 ;
        RECT 1.044 0.108 1.192 0.18 ;
        RECT 0.072 0.54 0.896 0.612 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V1 ;
        RECT 0.172 0.108 0.244 0.18 ;
        RECT 1.06 0.108 1.132 0.18 ;
      LAYER V0 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.396 0.54 0.468 0.612 ;
        RECT 0.824 0.54 0.896 0.612 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.612 0.396 0.872 0.468 ;
      LAYER M1 ;
        RECT 0.592 0.396 0.812 0.468 ;
      LAYER V1 ;
        RECT 0.612 0.396 0.684 0.468 ;
      LAYER V0 ;
        RECT 0.612 0.396 0.684 0.468 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 1.548 0.756 ;
      RECT 0.396 0.108 0.9 0.18 ;
  END
END AOI32x1_ASAP7_6t_fix

MACRO AOI32xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.328 0.396 0.596 0.468 ;
        RECT 0.328 0.54 0.548 0.612 ;
        RECT 0.328 0.108 0.476 0.18 ;
        RECT 0.328 0.108 0.4 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.54 1.028 0.612 ;
        RECT 0.792 0.252 1.028 0.324 ;
        RECT 0.792 0.252 0.864 0.612 ;
      LAYER V0 ;
        RECT 0.792 0.396 0.864 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.424 0.324 ;
        RECT 1.152 0.54 1.332 0.612 ;
        RECT 1.152 0.252 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.724 0.54 1.872 0.612 ;
        RECT 1.8 0.108 1.872 0.612 ;
        RECT 1.724 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 0.816 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.54 1.62 0.612 ;
        RECT 1.548 0.108 1.62 0.612 ;
        RECT 0.612 0.108 1.62 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.476 0.54 1.548 0.612 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 1.764 0.756 ;
  END
END AOI32xp33_ASAP7_6t_fix

MACRO AOI32xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32xp67_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.54 1.548 0.612 ;
        RECT 1.12 0.252 1.268 0.324 ;
        RECT 1.152 0.252 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.468 1.224 0.54 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.108 1.872 0.18 ;
        RECT 1.368 0.108 1.44 0.44 ;
      LAYER V0 ;
        RECT 1.368 0.34 1.44 0.412 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.684 1.872 0.756 ;
        RECT 1.8 0.252 1.872 0.756 ;
        RECT 1.54 0.252 1.872 0.324 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.46 ;
        RECT 0.288 0.252 1.008 0.324 ;
        RECT 0.288 0.252 0.36 0.44 ;
      LAYER V0 ;
        RECT 0.288 0.324 0.36 0.396 ;
        RECT 0.936 0.388 1.008 0.46 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.68 0.648 1.776 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.6 -0.048 0.696 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.152 0.108 1.144 0.18 ;
      LAYER M1 ;
        RECT 1.044 0.108 1.192 0.18 ;
        RECT 0.072 0.54 0.872 0.612 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V1 ;
        RECT 0.172 0.108 0.244 0.18 ;
        RECT 1.052 0.108 1.124 0.18 ;
      LAYER V0 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.396 0.54 0.468 0.612 ;
        RECT 0.78 0.54 0.852 0.612 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.268 0.396 1.06 0.468 ;
      LAYER M1 ;
        RECT 0.484 0.396 0.812 0.468 ;
      LAYER V1 ;
        RECT 0.612 0.396 0.684 0.468 ;
      LAYER V0 ;
        RECT 0.612 0.396 0.684 0.468 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 1.548 0.756 ;
      RECT 0.396 0.108 0.9 0.18 ;
  END
END AOI32xp67_ASAP7_6t_fix

MACRO AOI331xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI331xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.696 0.108 0.768 0.488 ;
        RECT 0.604 0.108 0.768 0.18 ;
      LAYER V0 ;
        RECT 0.696 0.396 0.768 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.296 0.576 0.584 ;
      LAYER V0 ;
        RECT 0.504 0.392 0.576 0.464 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.22 0.612 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.84 0.396 1.004 0.468 ;
        RECT 0.84 0.108 0.988 0.18 ;
        RECT 0.84 0.108 0.912 0.468 ;
      LAYER V0 ;
        RECT 0.912 0.396 0.984 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.104 0.396 1.268 0.468 ;
        RECT 1.104 0.312 1.176 0.468 ;
      LAYER V0 ;
        RECT 1.176 0.396 1.248 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.532 0.324 ;
        RECT 1.368 0.252 1.44 0.54 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.252 1.876 0.324 ;
        RECT 1.656 0.252 1.728 0.468 ;
      LAYER V0 ;
        RECT 1.656 0.396 1.728 0.468 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.108 1.764 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.524 0.532 1.596 0.704 ;
      RECT 0.396 0.684 1.332 0.756 ;
      RECT 0.972 0.54 1.18 0.612 ;
    LAYER M2 ;
      RECT 1.024 0.54 1.616 0.612 ;
    LAYER V1 ;
      RECT 1.524 0.54 1.596 0.612 ;
      RECT 1.044 0.54 1.116 0.612 ;
  END
END AOI331xp33_ASAP7_6t_fix

MACRO AOI332xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI332xp33_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.692 0.108 0.764 0.488 ;
        RECT 0.428 0.108 0.764 0.18 ;
      LAYER V0 ;
        RECT 0.692 0.396 0.764 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.244 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.292 0.18 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.108 1.136 0.18 ;
        RECT 0.86 0.396 1.008 0.468 ;
        RECT 0.86 0.108 0.936 0.468 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.252 1.72 0.324 ;
        RECT 1.132 0.396 1.368 0.468 ;
        RECT 1.296 0.252 1.368 0.468 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.588 0.54 1.808 0.612 ;
        RECT 1.736 0.396 1.808 0.612 ;
        RECT 1.492 0.396 1.808 0.468 ;
      LAYER V0 ;
        RECT 1.512 0.396 1.584 0.468 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.136 2.52 0.56 ;
      LAYER V0 ;
        RECT 2.448 0.396 2.52 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.844 0.252 2.204 0.324 ;
        RECT 1.908 0.54 2.056 0.612 ;
        RECT 1.984 0.252 2.056 0.612 ;
      LAYER V0 ;
        RECT 1.984 0.384 2.056 0.456 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 1.464 -0.048 1.992 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.156 0.54 2.376 0.612 ;
        RECT 2.304 0.108 2.376 0.612 ;
        RECT 1.26 0.108 2.376 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 2.156 0.54 2.228 0.612 ;
        RECT 2.304 0.252 2.376 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.908 0.756 ;
      RECT 0.836 0.54 0.908 0.756 ;
      RECT 0.836 0.54 1.376 0.612 ;
      RECT 1.044 0.684 2.412 0.756 ;
  END
END AOI332xp33_ASAP7_6t_fix

MACRO AOI333xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI333xp33_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.996 0.396 2.304 0.468 ;
        RECT 2.232 0.108 2.304 0.468 ;
        RECT 1.984 0.108 2.304 0.18 ;
      LAYER V0 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.836 0.396 1.028 0.468 ;
        RECT 0.836 0.396 0.908 0.544 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.432 ;
        RECT 0.928 0.252 1.224 0.324 ;
      LAYER V0 ;
        RECT 1.152 0.34 1.224 0.412 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.672 0.108 0.82 0.18 ;
        RECT 0.692 0.108 0.764 0.476 ;
      LAYER V0 ;
        RECT 0.692 0.384 0.764 0.456 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.256 0.576 0.472 ;
        RECT 0.428 0.256 0.576 0.328 ;
        RECT 0.428 0.108 0.5 0.328 ;
        RECT 0.072 0.108 0.5 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.4 0.576 0.472 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.288 0.324 ;
        RECT 0.072 0.252 0.144 0.62 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.124 0.684 2.308 0.756 ;
        RECT 2.124 0.54 2.196 0.756 ;
        RECT 1.712 0.54 2.196 0.612 ;
      LAYER V0 ;
        RECT 1.732 0.54 1.804 0.612 ;
        RECT 2.124 0.612 2.196 0.684 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.78 0.252 2.016 0.324 ;
      LAYER M1 ;
        RECT 1.8 0.252 1.948 0.324 ;
        RECT 1.8 0.252 1.872 0.44 ;
      LAYER V1 ;
        RECT 1.868 0.252 1.94 0.324 ;
      LAYER V0 ;
        RECT 1.8 0.348 1.872 0.42 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.54 0.396 1.872 0.468 ;
      LAYER M1 ;
        RECT 1.584 0.332 1.656 0.476 ;
      LAYER V1 ;
        RECT 1.584 0.396 1.656 0.468 ;
      LAYER V0 ;
        RECT 1.584 0.384 1.656 0.456 ;
    END
  END A3
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.156 0.252 1.54 0.324 ;
      LAYER M1 ;
        RECT 1.324 0.252 1.472 0.324 ;
        RECT 1.384 0.252 1.456 0.476 ;
      LAYER V1 ;
        RECT 1.384 0.252 1.456 0.324 ;
      LAYER V0 ;
        RECT 1.384 0.384 1.456 0.456 ;
    END
  END B3
  OBS
    LAYER M1 ;
      RECT 0.288 0.684 0.9 0.756 ;
      RECT 0.288 0.532 0.36 0.756 ;
      RECT 1.044 0.684 1.98 0.756 ;
      RECT 0.988 0.108 1.764 0.18 ;
      RECT 1.184 0.54 1.332 0.612 ;
    LAYER M2 ;
      RECT 0.268 0.54 1.332 0.612 ;
    LAYER V1 ;
      RECT 1.24 0.54 1.312 0.612 ;
      RECT 0.288 0.54 0.36 0.612 ;
  END
END AOI333xp33_ASAP7_6t_fix

MACRO AOI33x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33x1_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.372 0.756 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 1.116 0.468 ;
        RECT 0.36 0.54 0.66 0.612 ;
        RECT 0.36 0.252 0.66 0.324 ;
        RECT 0.36 0.252 0.432 0.612 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.396 1.76 0.468 ;
        RECT 1.508 0.54 1.656 0.612 ;
        RECT 1.584 0.396 1.656 0.612 ;
      LAYER V0 ;
        RECT 1.688 0.396 1.76 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.396 2.3 0.468 ;
        RECT 1.94 0.54 2.088 0.612 ;
        RECT 2.016 0.396 2.088 0.612 ;
      LAYER V0 ;
        RECT 2.204 0.396 2.276 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.252 2.52 0.44 ;
        RECT 2.232 0.252 2.52 0.324 ;
      LAYER V0 ;
        RECT 2.448 0.348 2.52 0.42 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.88 0.172 2.952 0.468 ;
      LAYER V0 ;
        RECT 2.88 0.396 2.952 0.468 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.752 0.54 2.824 0.684 ;
        RECT 2.296 0.54 2.824 0.612 ;
        RECT 2.664 0.108 2.736 0.612 ;
        RECT 1.672 0.108 2.736 0.18 ;
      LAYER V0 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.34 0.54 2.412 0.612 ;
        RECT 2.752 0.612 2.824 0.684 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.592 0.684 2.628 0.756 ;
      RECT 1.044 0.252 1.98 0.324 ;
      RECT 0.396 0.108 1.352 0.18 ;
  END
END AOI33x1_ASAP7_6t_fix

MACRO AOI33xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.288 0.18 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.108 0.576 0.42 ;
        RECT 0.412 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.348 0.576 0.42 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.604 0.54 0.768 0.612 ;
        RECT 0.696 0.136 0.768 0.612 ;
      LAYER V0 ;
        RECT 0.696 0.396 0.768 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.84 0.388 1.004 0.46 ;
        RECT 0.84 0.108 1.004 0.18 ;
        RECT 0.84 0.108 0.912 0.46 ;
      LAYER V0 ;
        RECT 0.912 0.388 0.984 0.46 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.104 0.396 1.268 0.468 ;
        RECT 1.104 0.24 1.176 0.468 ;
      LAYER V0 ;
        RECT 1.176 0.396 1.248 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.392 0.396 1.54 0.468 ;
        RECT 1.468 0.308 1.54 0.468 ;
      LAYER V0 ;
        RECT 1.392 0.396 1.464 0.468 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.684 1.684 0.756 ;
        RECT 1.612 0.108 1.684 0.756 ;
        RECT 1.004 0.54 1.684 0.612 ;
        RECT 1.26 0.108 1.684 0.18 ;
      LAYER V0 ;
        RECT 1.04 0.54 1.112 0.612 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.476 0.684 1.548 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 1.332 0.756 ;
  END
END AOI33xp33_ASAP7_6t_fix

MACRO ASYNC_DFFHx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ASYNC_DFFHx1_ASAP7_6t_fix 0 0 ;
  SIZE 5.832 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.36 0.756 ;
        RECT 0.288 0.488 0.36 0.756 ;
        RECT 0.072 0.108 0.276 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.508 0.36 0.58 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.408 1.152 0.48 ;
        RECT 0.936 0.252 1.008 0.48 ;
        RECT 0.648 0.252 1.008 0.324 ;
        RECT 0.648 0.252 0.72 0.612 ;
        RECT 0.5 0.684 0.648 0.756 ;
        RECT 0.576 0.54 0.648 0.756 ;
      LAYER V0 ;
        RECT 1.08 0.408 1.152 0.48 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.56 0.684 5.76 0.756 ;
        RECT 5.688 0.108 5.76 0.756 ;
        RECT 5.56 0.108 5.76 0.18 ;
      LAYER V0 ;
        RECT 5.58 0.684 5.652 0.756 ;
        RECT 5.58 0.108 5.652 0.18 ;
    END
  END QN
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.248 0.108 4.396 0.468 ;
        RECT 3.18 0.684 4.248 0.756 ;
        RECT 4.176 0.396 4.248 0.756 ;
        RECT 3.18 0.512 3.252 0.756 ;
        RECT 2.88 0.512 3.252 0.584 ;
        RECT 2.732 0.54 2.988 0.612 ;
      LAYER V0 ;
        RECT 2.796 0.54 2.868 0.612 ;
        RECT 3.096 0.512 3.168 0.584 ;
        RECT 4.176 0.516 4.248 0.588 ;
    END
  END SET
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 5.832 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 5.832 0.912 ;
        RECT 5.352 0.54 5.448 0.912 ;
        RECT 4.272 0.648 4.368 0.912 ;
        RECT 2.544 0.648 2.64 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.832 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 5.832 0.048 ;
        RECT 5.352 -0.048 5.448 0.324 ;
        RECT 4.704 -0.048 4.8 0.216 ;
        RECT 4.272 -0.048 4.368 0.216 ;
        RECT 2.976 -0.048 3.072 0.216 ;
        RECT 2.544 -0.048 2.64 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
    END
  END VSS
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.3 0.684 4.48 0.756 ;
      LAYER M1 ;
        RECT 4.38 0.684 4.536 0.756 ;
        RECT 4.464 0.516 4.536 0.756 ;
        RECT 2.3 0.684 2.488 0.756 ;
        RECT 2.416 0.496 2.488 0.756 ;
      LAYER V1 ;
        RECT 2.324 0.684 2.396 0.756 ;
        RECT 4.388 0.684 4.46 0.756 ;
      LAYER V0 ;
        RECT 2.416 0.516 2.488 0.588 ;
        RECT 4.464 0.516 4.536 0.588 ;
    END
  END RESET
  OBS
    LAYER M1 ;
      RECT 4.608 0.684 5.38 0.756 ;
      RECT 5.308 0.52 5.38 0.756 ;
      RECT 4.608 0.328 4.68 0.756 ;
      RECT 5.308 0.52 5.544 0.592 ;
      RECT 5.472 0.372 5.544 0.592 ;
      RECT 5 0.108 5.072 0.252 ;
      RECT 5 0.108 5.18 0.18 ;
      RECT 4.824 0.54 4.992 0.612 ;
      RECT 4.824 0.108 4.896 0.612 ;
      RECT 4.5 0.108 4.896 0.18 ;
      RECT 3.884 0.396 4.104 0.468 ;
      RECT 4.032 0.108 4.104 0.468 ;
      RECT 3.852 0.108 4.104 0.18 ;
      RECT 3.604 0.54 3.756 0.612 ;
      RECT 3.684 0.432 3.756 0.612 ;
      RECT 3.24 0.328 3.492 0.4 ;
      RECT 3.42 0.244 3.492 0.4 ;
      RECT 2.56 0.684 3.08 0.756 ;
      RECT 2.56 0.396 2.632 0.756 ;
      RECT 2.56 0.396 2.8 0.468 ;
      RECT 2.728 0.28 2.8 0.468 ;
      RECT 1.724 0.108 1.796 0.704 ;
      RECT 1.724 0.56 2.188 0.632 ;
      RECT 2.116 0.252 2.188 0.632 ;
      RECT 2.948 0.108 3.02 0.356 ;
      RECT 2.116 0.252 2.608 0.324 ;
      RECT 2.536 0.108 2.608 0.324 ;
      RECT 2.536 0.108 3.02 0.18 ;
      RECT 1.476 0.108 1.796 0.18 ;
      RECT 1.868 0.252 1.94 0.416 ;
      RECT 1.868 0.252 2.016 0.324 ;
      RECT 0.808 0.684 1.572 0.756 ;
      RECT 1.5 0.54 1.572 0.756 ;
      RECT 1.5 0.54 1.652 0.612 ;
      RECT 1.58 0.408 1.652 0.612 ;
      RECT 1.34 0.252 1.412 0.456 ;
      RECT 0.468 0.108 0.54 0.396 ;
      RECT 1.196 0.252 1.412 0.324 ;
      RECT 1.196 0.108 1.268 0.324 ;
      RECT 0.468 0.108 1.268 0.18 ;
      RECT 3.884 0.54 4.032 0.612 ;
      RECT 3.12 0.108 3.296 0.18 ;
      RECT 1.908 0.108 2.412 0.18 ;
    LAYER M2 ;
      RECT 3.128 0.108 5.172 0.18 ;
      RECT 3.872 0.54 4.984 0.612 ;
      RECT 2.568 0.396 3.984 0.468 ;
      RECT 1.572 0.54 3.732 0.612 ;
      RECT 1.332 0.252 3.54 0.324 ;
    LAYER V1 ;
      RECT 5.1 0.108 5.172 0.18 ;
      RECT 4.912 0.54 4.984 0.612 ;
      RECT 3.892 0.396 3.964 0.468 ;
      RECT 3.892 0.54 3.964 0.612 ;
      RECT 3.64 0.54 3.712 0.612 ;
      RECT 3.42 0.252 3.492 0.324 ;
      RECT 3.128 0.108 3.2 0.18 ;
      RECT 2.568 0.396 2.64 0.468 ;
      RECT 1.936 0.252 2.008 0.324 ;
      RECT 1.572 0.54 1.644 0.612 ;
      RECT 1.332 0.252 1.404 0.324 ;
  END
END ASYNC_DFFHx1_ASAP7_6t_fix

MACRO ASYNC_DFFHx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ASYNC_DFFHx2_ASAP7_6t_fix 0 0 ;
  SIZE 6.048 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.36 0.756 ;
        RECT 0.288 0.488 0.36 0.756 ;
        RECT 0.072 0.108 0.276 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.508 0.36 0.58 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.408 1.152 0.48 ;
        RECT 0.936 0.252 1.008 0.48 ;
        RECT 0.648 0.252 1.008 0.324 ;
        RECT 0.648 0.252 0.72 0.612 ;
        RECT 0.5 0.684 0.648 0.756 ;
        RECT 0.576 0.54 0.648 0.756 ;
      LAYER V0 ;
        RECT 1.08 0.408 1.152 0.48 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.56 0.684 5.904 0.756 ;
        RECT 5.832 0.108 5.904 0.756 ;
        RECT 5.56 0.108 5.904 0.18 ;
      LAYER V0 ;
        RECT 5.58 0.684 5.652 0.756 ;
        RECT 5.58 0.108 5.652 0.18 ;
    END
  END QN
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.248 0.18 4.396 0.468 ;
        RECT 3.18 0.684 4.248 0.756 ;
        RECT 4.176 0.396 4.248 0.756 ;
        RECT 3.18 0.512 3.252 0.756 ;
        RECT 2.88 0.512 3.252 0.584 ;
        RECT 2.732 0.54 2.988 0.612 ;
      LAYER V0 ;
        RECT 2.796 0.54 2.868 0.612 ;
        RECT 3.096 0.512 3.168 0.584 ;
        RECT 4.176 0.516 4.248 0.588 ;
    END
  END SET
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 6.048 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 6.048 0.912 ;
        RECT 5.784 0.54 5.88 0.912 ;
        RECT 5.352 0.54 5.448 0.912 ;
        RECT 4.272 0.648 4.368 0.912 ;
        RECT 2.544 0.648 2.64 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
        RECT 5.796 0.828 5.868 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.048 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 6.048 0.048 ;
        RECT 5.784 -0.048 5.88 0.324 ;
        RECT 5.352 -0.048 5.448 0.324 ;
        RECT 4.704 -0.048 4.8 0.216 ;
        RECT 4.272 -0.048 4.368 0.216 ;
        RECT 2.976 -0.048 3.072 0.216 ;
        RECT 2.544 -0.048 2.64 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
        RECT 5.796 -0.036 5.868 0.036 ;
    END
  END VSS
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.3 0.684 4.48 0.756 ;
      LAYER M1 ;
        RECT 4.38 0.684 4.536 0.756 ;
        RECT 4.464 0.516 4.536 0.756 ;
        RECT 2.3 0.684 2.488 0.756 ;
        RECT 2.416 0.496 2.488 0.756 ;
      LAYER V1 ;
        RECT 2.324 0.684 2.396 0.756 ;
        RECT 4.388 0.684 4.46 0.756 ;
      LAYER V0 ;
        RECT 2.416 0.516 2.488 0.588 ;
        RECT 4.464 0.516 4.536 0.588 ;
    END
  END RESET
  OBS
    LAYER M1 ;
      RECT 4.608 0.684 5.38 0.756 ;
      RECT 5.308 0.52 5.38 0.756 ;
      RECT 4.608 0.328 4.68 0.756 ;
      RECT 5.308 0.52 5.544 0.592 ;
      RECT 5.472 0.372 5.544 0.592 ;
      RECT 5 0.108 5.072 0.252 ;
      RECT 5 0.108 5.18 0.18 ;
      RECT 4.824 0.54 4.992 0.612 ;
      RECT 4.824 0.108 4.896 0.612 ;
      RECT 4.5 0.108 4.896 0.18 ;
      RECT 3.884 0.396 4.104 0.468 ;
      RECT 4.032 0.108 4.104 0.468 ;
      RECT 3.852 0.108 4.104 0.18 ;
      RECT 3.604 0.54 3.756 0.612 ;
      RECT 3.684 0.432 3.756 0.612 ;
      RECT 3.24 0.328 3.492 0.4 ;
      RECT 3.42 0.244 3.492 0.4 ;
      RECT 2.56 0.684 3.08 0.756 ;
      RECT 2.56 0.396 2.632 0.756 ;
      RECT 2.56 0.396 2.8 0.468 ;
      RECT 2.728 0.28 2.8 0.468 ;
      RECT 1.724 0.108 1.796 0.704 ;
      RECT 1.724 0.56 2.188 0.632 ;
      RECT 2.116 0.252 2.188 0.632 ;
      RECT 2.948 0.108 3.02 0.356 ;
      RECT 2.116 0.252 2.608 0.324 ;
      RECT 2.536 0.108 2.608 0.324 ;
      RECT 2.536 0.108 3.02 0.18 ;
      RECT 1.476 0.108 1.796 0.18 ;
      RECT 1.868 0.252 1.94 0.416 ;
      RECT 1.868 0.252 2.016 0.324 ;
      RECT 0.808 0.684 1.572 0.756 ;
      RECT 1.5 0.54 1.572 0.756 ;
      RECT 1.5 0.54 1.652 0.612 ;
      RECT 1.58 0.408 1.652 0.612 ;
      RECT 1.34 0.252 1.412 0.456 ;
      RECT 0.468 0.108 0.54 0.396 ;
      RECT 1.196 0.252 1.412 0.324 ;
      RECT 1.196 0.108 1.268 0.324 ;
      RECT 0.468 0.108 1.268 0.18 ;
      RECT 3.884 0.54 4.032 0.612 ;
      RECT 3.12 0.108 3.296 0.18 ;
      RECT 1.908 0.108 2.412 0.18 ;
    LAYER M2 ;
      RECT 3.128 0.108 5.172 0.18 ;
      RECT 3.872 0.54 4.984 0.612 ;
      RECT 2.568 0.396 3.984 0.468 ;
      RECT 1.572 0.54 3.732 0.612 ;
      RECT 1.332 0.252 3.54 0.324 ;
    LAYER V1 ;
      RECT 5.1 0.108 5.172 0.18 ;
      RECT 4.912 0.54 4.984 0.612 ;
      RECT 3.892 0.396 3.964 0.468 ;
      RECT 3.892 0.54 3.964 0.612 ;
      RECT 3.64 0.54 3.712 0.612 ;
      RECT 3.42 0.252 3.492 0.324 ;
      RECT 3.128 0.108 3.2 0.18 ;
      RECT 2.568 0.396 2.64 0.468 ;
      RECT 1.936 0.252 2.008 0.324 ;
      RECT 1.572 0.54 1.644 0.612 ;
      RECT 1.332 0.252 1.404 0.324 ;
  END
END ASYNC_DFFHx2_ASAP7_6t_fix

MACRO BUFx10_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx10_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.684 2.736 0.756 ;
        RECT 2.664 0.108 2.736 0.756 ;
        RECT 0.796 0.108 2.736 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.576 0.756 ;
      RECT 0.504 0.108 0.576 0.756 ;
      RECT 0.504 0.396 0.792 0.468 ;
      RECT 0.396 0.108 0.576 0.18 ;
  END
END BUFx10_ASAP7_6t_fix

MACRO BUFx12_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.684 3.168 0.756 ;
        RECT 3.096 0.108 3.168 0.756 ;
        RECT 0.796 0.108 3.168 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 0.576 0.756 ;
      RECT 0.504 0.108 0.576 0.756 ;
      RECT 0.504 0.396 0.792 0.468 ;
      RECT 0.376 0.108 0.576 0.18 ;
  END
END BUFx12_ASAP7_6t_fix

MACRO BUFx12f_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx12f_ASAP7_6t_fix 0 0 ;
  SIZE 3.888 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.888 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.888 0.912 ;
        RECT 3.624 0.54 3.72 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.888 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.888 0.048 ;
        RECT 3.624 -0.048 3.72 0.324 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 3.824 0.756 ;
        RECT 1.24 0.108 3.824 0.18 ;
        RECT 3.744 0.108 3.816 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
        RECT 3.42 0.684 3.492 0.756 ;
        RECT 3.42 0.108 3.492 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 1.116 0.756 ;
      RECT 1.044 0.108 1.116 0.756 ;
      RECT 1.044 0.396 1.244 0.468 ;
      RECT 0.376 0.108 1.116 0.18 ;
  END
END BUFx12f_ASAP7_6t_fix

MACRO BUFx16f_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx16f_ASAP7_6t_fix 0 0 ;
  SIZE 4.752 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.752 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.752 0.912 ;
        RECT 4.488 0.54 4.584 0.912 ;
        RECT 4.056 0.54 4.152 0.912 ;
        RECT 3.624 0.54 3.72 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.752 0.048 ;
        RECT 4.488 -0.048 4.584 0.324 ;
        RECT 4.056 -0.048 4.152 0.324 ;
        RECT 3.624 -0.048 3.72 0.324 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 4.68 0.756 ;
        RECT 4.608 0.108 4.68 0.756 ;
        RECT 1.24 0.108 4.68 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
        RECT 3.42 0.684 3.492 0.756 ;
        RECT 3.42 0.108 3.492 0.18 ;
        RECT 3.852 0.684 3.924 0.756 ;
        RECT 3.852 0.108 3.924 0.18 ;
        RECT 4.284 0.684 4.356 0.756 ;
        RECT 4.284 0.108 4.356 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 1.008 0.756 ;
      RECT 0.936 0.108 1.008 0.756 ;
      RECT 0.936 0.396 1.224 0.468 ;
      RECT 0.376 0.108 1.008 0.18 ;
  END
END BUFx16f_ASAP7_6t_fix

MACRO BUFx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx1_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.404 0.468 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.288 0.396 0.36 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.684 0.792 0.756 ;
        RECT 0.72 0.108 0.792 0.756 ;
        RECT 0.644 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.084 0.54 0.576 0.612 ;
      RECT 0.504 0.28 0.576 0.612 ;
  END
END BUFx1_ASAP7_6t_fix

MACRO BUFx24_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx24_ASAP7_6t_fix 0 0 ;
  SIZE 6.48 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 6.48 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 6.48 0.912 ;
        RECT 6.216 0.54 6.312 0.912 ;
        RECT 5.784 0.54 5.88 0.912 ;
        RECT 5.352 0.54 5.448 0.912 ;
        RECT 4.92 0.54 5.016 0.912 ;
        RECT 4.488 0.54 4.584 0.912 ;
        RECT 4.056 0.54 4.152 0.912 ;
        RECT 3.624 0.54 3.72 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
        RECT 5.796 0.828 5.868 0.9 ;
        RECT 6.012 0.828 6.084 0.9 ;
        RECT 6.228 0.828 6.3 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.48 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 6.48 0.048 ;
        RECT 6.216 -0.048 6.312 0.324 ;
        RECT 5.784 -0.048 5.88 0.324 ;
        RECT 5.352 -0.048 5.448 0.324 ;
        RECT 4.92 -0.048 5.016 0.324 ;
        RECT 4.488 -0.048 4.584 0.324 ;
        RECT 4.056 -0.048 4.152 0.324 ;
        RECT 3.624 -0.048 3.72 0.324 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
        RECT 5.796 -0.036 5.868 0.036 ;
        RECT 6.012 -0.036 6.084 0.036 ;
        RECT 6.228 -0.036 6.3 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 6.408 0.756 ;
        RECT 6.336 0.108 6.408 0.756 ;
        RECT 1.24 0.108 6.408 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
        RECT 3.42 0.684 3.492 0.756 ;
        RECT 3.42 0.108 3.492 0.18 ;
        RECT 3.852 0.684 3.924 0.756 ;
        RECT 3.852 0.108 3.924 0.18 ;
        RECT 4.284 0.684 4.356 0.756 ;
        RECT 4.284 0.108 4.356 0.18 ;
        RECT 4.716 0.684 4.788 0.756 ;
        RECT 4.716 0.108 4.788 0.18 ;
        RECT 5.148 0.684 5.22 0.756 ;
        RECT 5.148 0.108 5.22 0.18 ;
        RECT 5.58 0.684 5.652 0.756 ;
        RECT 5.58 0.108 5.652 0.18 ;
        RECT 6.012 0.684 6.084 0.756 ;
        RECT 6.012 0.108 6.084 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 1.008 0.756 ;
      RECT 0.936 0.108 1.008 0.756 ;
      RECT 0.936 0.396 1.224 0.468 ;
      RECT 0.376 0.108 1.008 0.18 ;
  END
END BUFx24_ASAP7_6t_fix

MACRO BUFx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.612 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.228 0.268 0.3 0.596 ;
      RECT 0.228 0.396 0.792 0.468 ;
  END
END BUFx2_ASAP7_6t_fix

MACRO BUFx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 0.592 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.228 0.268 0.3 0.596 ;
      RECT 0.228 0.396 0.576 0.468 ;
  END
END BUFx3_ASAP7_6t_fix

MACRO BUFx4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 0.612 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.228 0.268 0.3 0.596 ;
      RECT 0.228 0.396 0.576 0.468 ;
  END
END BUFx4_ASAP7_6t_fix

MACRO BUFx4f_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4f_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.608 0.212 0.756 ;
        RECT 0.064 0.108 0.212 0.256 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.684 1.664 0.756 ;
        RECT 0.796 0.108 1.664 0.18 ;
        RECT 1.584 0.108 1.656 0.756 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.576 0.756 ;
      RECT 0.504 0.108 0.576 0.756 ;
      RECT 0.504 0.396 0.792 0.468 ;
      RECT 0.396 0.108 0.576 0.18 ;
  END
END BUFx4f_ASAP7_6t_fix

MACRO BUFx5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx5_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 1.548 0.756 ;
        RECT 0.612 0.108 1.548 0.18 ;
        RECT 1.368 0.108 1.44 0.756 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.228 0.268 0.3 0.596 ;
      RECT 0.228 0.396 0.576 0.468 ;
  END
END BUFx5_ASAP7_6t_fix

MACRO BUFx6f_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx6f_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.328 0.468 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.236 0.396 0.308 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.684 2.088 0.756 ;
        RECT 2.016 0.108 2.088 0.756 ;
        RECT 0.808 0.108 2.088 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.576 0.756 ;
      RECT 0.504 0.108 0.576 0.756 ;
      RECT 0.504 0.396 0.792 0.468 ;
      RECT 0.396 0.108 0.576 0.18 ;
  END
END BUFx6f_ASAP7_6t_fix

MACRO BUFx8_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 2.528 0.756 ;
        RECT 0.828 0.108 2.528 0.18 ;
        RECT 2.448 0.108 2.52 0.756 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.576 0.756 ;
      RECT 0.504 0.108 0.576 0.756 ;
      RECT 0.504 0.396 0.792 0.468 ;
      RECT 0.396 0.108 0.576 0.18 ;
  END
END BUFx8_ASAP7_6t_fix

MACRO BUFxp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFxp33_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 0.8 0.756 ;
        RECT 0.592 0.108 0.8 0.18 ;
        RECT 0.72 0.108 0.792 0.756 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.228 0.268 0.3 0.596 ;
      RECT 0.228 0.396 0.576 0.468 ;
  END
END BUFxp33_ASAP7_6t_fix

MACRO BUFxp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFxp67_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 0.8 0.756 ;
        RECT 0.592 0.108 0.8 0.18 ;
        RECT 0.72 0.108 0.792 0.756 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.228 0.268 0.3 0.596 ;
      RECT 0.228 0.396 0.596 0.468 ;
  END
END BUFxp67_ASAP7_6t_fix

MACRO DECAPx10_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx10_ASAP7_6t_fix 0 0 ;
  SIZE 4.752 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.752 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.752 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.752 0.048 ;
        RECT 4.272 -0.048 4.368 0.324 ;
        RECT 3.84 -0.048 3.936 0.324 ;
        RECT 3.408 -0.048 3.504 0.324 ;
        RECT 2.976 -0.048 3.072 0.324 ;
        RECT 2.544 -0.048 2.64 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.232 0.18 2.304 0.488 ;
      RECT 2.232 0.18 4.592 0.252 ;
      RECT 0.16 0.612 2.52 0.684 ;
      RECT 2.448 0.376 2.52 0.684 ;
  END
END DECAPx10_ASAP7_6t_fix

MACRO DECAPx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx1_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.376 0.612 0.576 0.684 ;
      RECT 0.504 0.42 0.576 0.684 ;
      RECT 0.288 0.18 0.36 0.444 ;
      RECT 0.288 0.18 0.488 0.252 ;
  END
END DECAPx1_ASAP7_6t_fix

MACRO DECAPx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx2_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.504 0.18 0.576 0.444 ;
      RECT 0.504 0.18 1.136 0.252 ;
      RECT 0.16 0.612 0.792 0.684 ;
      RECT 0.72 0.376 0.792 0.684 ;
  END
END DECAPx2_ASAP7_6t_fix

MACRO DECAPx4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx4_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.936 0.18 1.008 0.488 ;
      RECT 0.936 0.18 2 0.252 ;
      RECT 0.16 0.612 1.224 0.684 ;
      RECT 1.152 0.376 1.224 0.684 ;
  END
END DECAPx4_ASAP7_6t_fix

MACRO DECAPx6_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAPx6_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 2.544 -0.048 2.64 0.324 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.368 0.18 1.44 0.488 ;
      RECT 1.368 0.18 2.864 0.252 ;
      RECT 0.16 0.612 1.656 0.684 ;
      RECT 1.584 0.376 1.656 0.684 ;
  END
END DECAPx6_ASAP7_6t_fix

MACRO DFFHQNx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1_ASAP7_6t_fix 0 0 ;
  SIZE 4.752 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.684 1.008 0.756 ;
        RECT 0.936 0.252 1.008 0.756 ;
        RECT 0.86 0.252 1.008 0.324 ;
      LAYER V0 ;
        RECT 0.936 0.324 1.008 0.396 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.528 0.684 4.68 0.756 ;
        RECT 4.608 0.108 4.68 0.756 ;
        RECT 4.528 0.108 4.68 0.18 ;
      LAYER V0 ;
        RECT 4.608 0.396 4.68 0.468 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.216 0.144 0.288 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.752 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.752 0.912 ;
        RECT 4.488 0.54 4.584 0.912 ;
        RECT 3.408 0.648 3.504 0.912 ;
        RECT 1.896 0.648 1.992 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.56 0.828 2.632 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.64 0.828 3.712 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.752 0.048 ;
        RECT 4.488 -0.048 4.584 0.324 ;
        RECT 3.408 -0.048 3.504 0.216 ;
        RECT 1.896 -0.048 1.992 0.216 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.852 0.684 4.392 0.756 ;
      RECT 4.32 0.108 4.392 0.756 ;
      RECT 3.312 0.108 3.384 0.356 ;
      RECT 3.312 0.108 4.392 0.18 ;
      RECT 3.096 0.54 3.54 0.612 ;
      RECT 3.468 0.272 3.54 0.612 ;
      RECT 2.664 0.324 2.736 0.58 ;
      RECT 3.096 0.324 3.168 0.612 ;
      RECT 4.176 0.272 4.248 0.488 ;
      RECT 1.152 0.324 1.224 0.472 ;
      RECT 1.152 0.324 3.168 0.396 ;
      RECT 3.468 0.272 4.248 0.344 ;
      RECT 1.36 0.684 3.728 0.756 ;
      RECT 3.656 0.416 3.728 0.756 ;
      RECT 2.88 0.508 2.952 0.756 ;
      RECT 2.232 0.52 2.304 0.756 ;
      RECT 1.36 0.576 1.432 0.756 ;
      RECT 3.656 0.416 4.032 0.488 ;
      RECT 0.288 0.252 0.36 0.484 ;
      RECT 0.288 0.252 0.468 0.324 ;
      RECT 0.396 0.108 0.468 0.324 ;
      RECT 0.396 0.108 2.844 0.18 ;
      RECT 1.596 0.52 2.088 0.592 ;
  END
END DFFHQNx1_ASAP7_6t_fix

MACRO DFFHQNx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2_ASAP7_6t_fix 0 0 ;
  SIZE 4.968 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.508 1.224 0.58 ;
        RECT 0.936 0.252 1.224 0.324 ;
        RECT 0.936 0.252 1.008 0.58 ;
        RECT 0.592 0.684 0.864 0.756 ;
        RECT 0.792 0.508 0.864 0.756 ;
      LAYER V0 ;
        RECT 1.152 0.508 1.224 0.58 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.748 0.684 4.896 0.756 ;
        RECT 4.824 0.108 4.896 0.756 ;
        RECT 4.748 0.108 4.896 0.18 ;
      LAYER V0 ;
        RECT 4.824 0.396 4.896 0.468 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.468 0.756 ;
        RECT 0.072 0.108 0.468 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.968 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.968 0.912 ;
        RECT 4.704 0.54 4.8 0.912 ;
        RECT 3.624 0.648 3.72 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.776 0.828 2.848 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.856 0.828 3.928 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.968 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.968 0.048 ;
        RECT 4.704 -0.048 4.8 0.324 ;
        RECT 3.624 -0.048 3.72 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.248 -0.048 1.344 0.216 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.068 0.684 4.608 0.756 ;
      RECT 4.536 0.108 4.608 0.756 ;
      RECT 3.528 0.108 3.6 0.356 ;
      RECT 3.528 0.108 4.608 0.18 ;
      RECT 1.044 0.684 1.44 0.756 ;
      RECT 1.368 0.324 1.44 0.756 ;
      RECT 3.312 0.54 3.756 0.612 ;
      RECT 3.684 0.272 3.756 0.612 ;
      RECT 2.88 0.324 2.952 0.58 ;
      RECT 3.312 0.324 3.384 0.612 ;
      RECT 4.392 0.272 4.464 0.488 ;
      RECT 1.368 0.324 3.384 0.396 ;
      RECT 3.684 0.272 4.464 0.344 ;
      RECT 1.576 0.684 3.944 0.756 ;
      RECT 3.872 0.416 3.944 0.756 ;
      RECT 3.096 0.508 3.168 0.756 ;
      RECT 2.448 0.52 2.52 0.756 ;
      RECT 1.576 0.576 1.648 0.756 ;
      RECT 3.872 0.416 4.248 0.488 ;
      RECT 0.504 0.392 0.684 0.464 ;
      RECT 0.612 0.108 0.684 0.464 ;
      RECT 0.612 0.108 3.06 0.18 ;
      RECT 1.812 0.52 2.304 0.592 ;
  END
END DFFHQNx2_ASAP7_6t_fix

MACRO DFFHQNx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3_ASAP7_6t_fix 0 0 ;
  SIZE 5.184 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.508 1.44 0.58 ;
        RECT 1.152 0.252 1.44 0.324 ;
        RECT 1.152 0.252 1.224 0.58 ;
        RECT 0.808 0.684 1.08 0.756 ;
        RECT 1.008 0.508 1.08 0.756 ;
      LAYER V0 ;
        RECT 1.368 0.508 1.44 0.58 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.96 0.684 5.112 0.756 ;
        RECT 5.04 0.108 5.112 0.756 ;
        RECT 4.96 0.108 5.112 0.18 ;
      LAYER V0 ;
        RECT 5.04 0.396 5.112 0.468 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.684 0.756 ;
        RECT 0.072 0.108 0.684 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 5.184 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 5.184 0.912 ;
        RECT 4.92 0.54 5.016 0.912 ;
        RECT 3.84 0.648 3.936 0.912 ;
        RECT 2.328 0.648 2.424 0.912 ;
        RECT 1.464 0.648 1.56 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.992 0.828 3.064 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.072 0.828 4.144 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.184 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 5.184 0.048 ;
        RECT 4.92 -0.048 5.016 0.324 ;
        RECT 3.84 -0.048 3.936 0.216 ;
        RECT 2.328 -0.048 2.424 0.216 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.284 0.684 4.824 0.756 ;
      RECT 4.752 0.108 4.824 0.756 ;
      RECT 3.744 0.108 3.816 0.356 ;
      RECT 3.744 0.108 4.824 0.18 ;
      RECT 1.26 0.684 1.656 0.756 ;
      RECT 1.584 0.324 1.656 0.756 ;
      RECT 3.528 0.54 3.972 0.612 ;
      RECT 3.9 0.272 3.972 0.612 ;
      RECT 3.096 0.324 3.168 0.58 ;
      RECT 3.528 0.324 3.6 0.612 ;
      RECT 4.608 0.272 4.68 0.488 ;
      RECT 1.584 0.324 3.6 0.396 ;
      RECT 3.9 0.272 4.68 0.344 ;
      RECT 1.792 0.684 4.16 0.756 ;
      RECT 4.088 0.416 4.16 0.756 ;
      RECT 3.312 0.508 3.384 0.756 ;
      RECT 2.664 0.52 2.736 0.756 ;
      RECT 1.792 0.576 1.864 0.756 ;
      RECT 4.088 0.416 4.464 0.488 ;
      RECT 0.72 0.392 0.9 0.464 ;
      RECT 0.828 0.108 0.9 0.464 ;
      RECT 0.828 0.108 3.276 0.18 ;
      RECT 2.028 0.52 2.52 0.592 ;
  END
END DFFHQNx3_ASAP7_6t_fix

MACRO DFFHQx4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQx4_ASAP7_6t_fix 0 0 ;
  SIZE 5.832 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.508 2.088 0.58 ;
        RECT 1.8 0.252 2.088 0.324 ;
        RECT 1.8 0.252 1.872 0.58 ;
        RECT 1.456 0.684 1.728 0.756 ;
        RECT 1.656 0.508 1.728 0.756 ;
      LAYER V0 ;
        RECT 2.016 0.508 2.088 0.58 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.608 0.684 5.76 0.756 ;
        RECT 5.688 0.108 5.76 0.756 ;
        RECT 5.608 0.108 5.76 0.18 ;
      LAYER V0 ;
        RECT 5.688 0.396 5.76 0.468 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.9 0.756 ;
        RECT 0.072 0.108 0.9 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 5.832 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 5.832 0.912 ;
        RECT 5.568 0.54 5.664 0.912 ;
        RECT 4.488 0.648 4.584 0.912 ;
        RECT 2.976 0.648 3.072 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.64 0.828 3.712 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.72 0.828 4.792 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.832 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 5.832 0.048 ;
        RECT 5.568 -0.048 5.664 0.324 ;
        RECT 4.488 -0.048 4.584 0.216 ;
        RECT 2.976 -0.048 3.072 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.932 0.684 5.472 0.756 ;
      RECT 5.4 0.108 5.472 0.756 ;
      RECT 4.392 0.108 4.464 0.356 ;
      RECT 4.392 0.108 5.472 0.18 ;
      RECT 1.908 0.684 2.304 0.756 ;
      RECT 2.232 0.324 2.304 0.756 ;
      RECT 4.176 0.54 4.62 0.612 ;
      RECT 4.548 0.272 4.62 0.612 ;
      RECT 3.744 0.324 3.816 0.58 ;
      RECT 4.176 0.324 4.248 0.612 ;
      RECT 5.256 0.272 5.328 0.488 ;
      RECT 2.232 0.324 4.248 0.396 ;
      RECT 4.548 0.272 5.328 0.344 ;
      RECT 2.44 0.684 4.808 0.756 ;
      RECT 4.736 0.416 4.808 0.756 ;
      RECT 3.96 0.508 4.032 0.756 ;
      RECT 3.312 0.52 3.384 0.756 ;
      RECT 2.44 0.576 2.512 0.756 ;
      RECT 4.736 0.416 5.112 0.488 ;
      RECT 1.368 0.392 1.548 0.464 ;
      RECT 1.476 0.108 1.548 0.464 ;
      RECT 1.476 0.108 3.924 0.18 ;
      RECT 1.044 0.684 1.332 0.756 ;
      RECT 1.044 0.108 1.116 0.756 ;
      RECT 0.72 0.392 1.116 0.464 ;
      RECT 1.044 0.108 1.332 0.18 ;
      RECT 2.676 0.52 3.168 0.592 ;
  END
END DFFHQx4_ASAP7_6t_fix

MACRO DFFLQNx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx1_ASAP7_6t_fix 0 0 ;
  SIZE 4.32 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.584 0.756 ;
        RECT 0.072 0.252 0.58 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.464 0.36 0.536 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.712 0.684 1.156 0.756 ;
        RECT 1.084 0.352 1.156 0.756 ;
      LAYER V0 ;
        RECT 1.084 0.392 1.156 0.464 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.684 4.248 0.756 ;
        RECT 4.176 0.108 4.248 0.756 ;
        RECT 4.048 0.108 4.248 0.18 ;
      LAYER V0 ;
        RECT 4.068 0.684 4.14 0.756 ;
        RECT 4.068 0.108 4.14 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.32 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.32 0.912 ;
        RECT 3.84 0.54 3.936 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.32 0.048 ;
        RECT 3.84 -0.048 3.936 0.324 ;
        RECT 3.192 -0.048 3.288 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.88 0.108 2.952 0.72 ;
      RECT 2.88 0.508 3.6 0.58 ;
      RECT 3.528 0.396 3.6 0.58 ;
      RECT 3.312 0.396 3.384 0.58 ;
      RECT 3.528 0.396 4.032 0.468 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 3.096 0.108 3.168 0.364 ;
      RECT 3.096 0.108 3.492 0.18 ;
      RECT 2.008 0.656 2.592 0.728 ;
      RECT 2.52 0.252 2.592 0.728 ;
      RECT 2.008 0.5 2.08 0.728 ;
      RECT 2.34 0.252 2.592 0.324 ;
      RECT 2.34 0.156 2.412 0.324 ;
      RECT 2.16 0.512 2.324 0.584 ;
      RECT 2.16 0.328 2.232 0.584 ;
      RECT 2.088 0.108 2.16 0.4 ;
      RECT 1.584 0.108 2.16 0.18 ;
      RECT 1.8 0.252 1.872 0.628 ;
      RECT 1.74 0.348 1.964 0.42 ;
      RECT 1.74 0.252 1.888 0.42 ;
      RECT 1.228 0.684 1.548 0.756 ;
      RECT 1.228 0.108 1.3 0.756 ;
      RECT 1.112 0.108 1.3 0.18 ;
      RECT 0.484 0.396 0.792 0.468 ;
      RECT 0.72 0.108 0.792 0.468 ;
      RECT 0.18 0.108 0.792 0.18 ;
      RECT 2.664 0.376 2.736 0.58 ;
      RECT 1.58 0.368 1.652 0.552 ;
      RECT 1.372 0.232 1.444 0.54 ;
      RECT 0.864 0.332 0.936 0.488 ;
    LAYER M2 ;
      RECT 0.844 0.396 2.756 0.468 ;
      RECT 0.7 0.252 1.896 0.324 ;
      RECT 1.12 0.108 1.76 0.18 ;
    LAYER V1 ;
      RECT 2.664 0.396 2.736 0.468 ;
      RECT 1.804 0.252 1.876 0.324 ;
      RECT 1.668 0.108 1.74 0.18 ;
      RECT 1.58 0.396 1.652 0.468 ;
      RECT 1.372 0.252 1.444 0.324 ;
      RECT 1.12 0.108 1.192 0.18 ;
      RECT 0.864 0.396 0.936 0.468 ;
      RECT 0.72 0.252 0.792 0.324 ;
  END
END DFFLQNx1_ASAP7_6t_fix

MACRO DFFLQNx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx2_ASAP7_6t_fix 0 0 ;
  SIZE 4.536 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.584 0.756 ;
        RECT 0.072 0.252 0.58 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.464 0.36 0.536 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.712 0.684 1.156 0.756 ;
        RECT 1.084 0.352 1.156 0.756 ;
      LAYER V0 ;
        RECT 1.084 0.392 1.156 0.464 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.684 4.464 0.756 ;
        RECT 4.392 0.108 4.464 0.756 ;
        RECT 4.048 0.108 4.464 0.18 ;
      LAYER V0 ;
        RECT 4.068 0.684 4.14 0.756 ;
        RECT 4.068 0.108 4.14 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.536 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.536 0.912 ;
        RECT 4.272 0.54 4.368 0.912 ;
        RECT 3.84 0.54 3.936 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.536 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.536 0.048 ;
        RECT 4.272 -0.048 4.368 0.324 ;
        RECT 3.84 -0.048 3.936 0.324 ;
        RECT 3.192 -0.048 3.288 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.88 0.108 2.952 0.72 ;
      RECT 2.88 0.508 3.6 0.58 ;
      RECT 3.528 0.396 3.6 0.58 ;
      RECT 3.312 0.396 3.384 0.58 ;
      RECT 3.528 0.396 4.032 0.468 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 3.096 0.108 3.168 0.364 ;
      RECT 3.096 0.108 3.492 0.18 ;
      RECT 2.008 0.656 2.592 0.728 ;
      RECT 2.52 0.252 2.592 0.728 ;
      RECT 2.008 0.5 2.08 0.728 ;
      RECT 2.34 0.252 2.592 0.324 ;
      RECT 2.34 0.156 2.412 0.324 ;
      RECT 2.16 0.512 2.324 0.584 ;
      RECT 2.16 0.328 2.232 0.584 ;
      RECT 2.088 0.108 2.16 0.4 ;
      RECT 1.584 0.108 2.16 0.18 ;
      RECT 1.8 0.252 1.872 0.628 ;
      RECT 1.74 0.348 1.964 0.42 ;
      RECT 1.74 0.252 1.888 0.42 ;
      RECT 1.228 0.684 1.548 0.756 ;
      RECT 1.228 0.108 1.3 0.756 ;
      RECT 1.112 0.108 1.3 0.18 ;
      RECT 0.484 0.396 0.792 0.468 ;
      RECT 0.72 0.108 0.792 0.468 ;
      RECT 0.18 0.108 0.792 0.18 ;
      RECT 2.664 0.376 2.736 0.58 ;
      RECT 1.58 0.368 1.652 0.552 ;
      RECT 1.372 0.232 1.444 0.54 ;
      RECT 0.864 0.332 0.936 0.488 ;
    LAYER M2 ;
      RECT 0.844 0.396 2.756 0.468 ;
      RECT 0.7 0.252 1.896 0.324 ;
      RECT 1.12 0.108 1.76 0.18 ;
    LAYER V1 ;
      RECT 2.664 0.396 2.736 0.468 ;
      RECT 1.804 0.252 1.876 0.324 ;
      RECT 1.668 0.108 1.74 0.18 ;
      RECT 1.58 0.396 1.652 0.468 ;
      RECT 1.372 0.252 1.444 0.324 ;
      RECT 1.12 0.108 1.192 0.18 ;
      RECT 0.864 0.396 0.936 0.468 ;
      RECT 0.72 0.252 0.792 0.324 ;
  END
END DFFLQNx2_ASAP7_6t_fix

MACRO DFFLQNx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQNx3_ASAP7_6t_fix 0 0 ;
  SIZE 4.752 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.584 0.756 ;
        RECT 0.072 0.252 0.58 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.464 0.36 0.536 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.712 0.684 1.156 0.756 ;
        RECT 1.084 0.352 1.156 0.756 ;
      LAYER V0 ;
        RECT 1.084 0.392 1.156 0.464 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.684 4.68 0.756 ;
        RECT 4.608 0.108 4.68 0.756 ;
        RECT 4.048 0.108 4.68 0.18 ;
      LAYER V0 ;
        RECT 4.068 0.684 4.14 0.756 ;
        RECT 4.068 0.108 4.14 0.18 ;
        RECT 4.5 0.684 4.572 0.756 ;
        RECT 4.5 0.108 4.572 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.752 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.752 0.912 ;
        RECT 4.272 0.54 4.368 0.912 ;
        RECT 3.84 0.54 3.936 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.752 0.048 ;
        RECT 4.272 -0.048 4.368 0.324 ;
        RECT 3.84 -0.048 3.936 0.324 ;
        RECT 3.192 -0.048 3.288 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.88 0.108 2.952 0.72 ;
      RECT 2.88 0.508 3.6 0.58 ;
      RECT 3.528 0.396 3.6 0.58 ;
      RECT 3.312 0.396 3.384 0.58 ;
      RECT 3.528 0.396 4.032 0.468 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 3.096 0.108 3.168 0.364 ;
      RECT 3.096 0.108 3.492 0.18 ;
      RECT 2.008 0.656 2.592 0.728 ;
      RECT 2.52 0.252 2.592 0.728 ;
      RECT 2.008 0.5 2.08 0.728 ;
      RECT 2.34 0.252 2.592 0.324 ;
      RECT 2.34 0.156 2.412 0.324 ;
      RECT 2.16 0.512 2.324 0.584 ;
      RECT 2.16 0.328 2.232 0.584 ;
      RECT 2.088 0.108 2.16 0.4 ;
      RECT 1.584 0.108 2.16 0.18 ;
      RECT 1.8 0.252 1.872 0.628 ;
      RECT 1.74 0.348 1.964 0.42 ;
      RECT 1.74 0.252 1.888 0.42 ;
      RECT 1.228 0.684 1.548 0.756 ;
      RECT 1.228 0.108 1.3 0.756 ;
      RECT 1.112 0.108 1.3 0.18 ;
      RECT 0.484 0.396 0.792 0.468 ;
      RECT 0.72 0.108 0.792 0.468 ;
      RECT 0.18 0.108 0.792 0.18 ;
      RECT 2.664 0.376 2.736 0.58 ;
      RECT 1.58 0.368 1.652 0.552 ;
      RECT 1.372 0.232 1.444 0.54 ;
      RECT 0.864 0.332 0.936 0.488 ;
    LAYER M2 ;
      RECT 0.844 0.396 2.756 0.468 ;
      RECT 0.7 0.252 1.896 0.324 ;
      RECT 1.12 0.108 1.76 0.18 ;
    LAYER V1 ;
      RECT 2.664 0.396 2.736 0.468 ;
      RECT 1.804 0.252 1.876 0.324 ;
      RECT 1.668 0.108 1.74 0.18 ;
      RECT 1.58 0.396 1.652 0.468 ;
      RECT 1.372 0.252 1.444 0.324 ;
      RECT 1.12 0.108 1.192 0.18 ;
      RECT 0.864 0.396 0.936 0.468 ;
      RECT 0.72 0.252 0.792 0.324 ;
  END
END DFFLQNx3_ASAP7_6t_fix

MACRO DFFLQx4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQx4_ASAP7_6t_fix 0 0 ;
  SIZE 5.4 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.584 0.756 ;
        RECT 0.072 0.252 0.58 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.464 0.36 0.536 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.712 0.684 1.156 0.756 ;
        RECT 1.084 0.352 1.156 0.756 ;
      LAYER V0 ;
        RECT 1.084 0.392 1.156 0.464 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5 0.684 5.328 0.756 ;
        RECT 5.256 0.108 5.328 0.756 ;
        RECT 4.5 0.108 5.328 0.18 ;
        RECT 4.5 0.592 4.572 0.756 ;
        RECT 4.5 0.108 4.572 0.272 ;
      LAYER V0 ;
        RECT 4.5 0.612 4.572 0.684 ;
        RECT 4.5 0.18 4.572 0.252 ;
        RECT 4.932 0.684 5.004 0.756 ;
        RECT 4.932 0.108 5.004 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 5.4 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 5.4 0.912 ;
        RECT 5.136 0.54 5.232 0.912 ;
        RECT 4.704 0.54 4.8 0.912 ;
        RECT 4.272 0.54 4.368 0.912 ;
        RECT 3.84 0.54 3.936 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 5.4 0.048 ;
        RECT 5.136 -0.048 5.232 0.324 ;
        RECT 4.704 -0.048 4.8 0.324 ;
        RECT 4.272 -0.048 4.368 0.324 ;
        RECT 3.84 -0.048 3.936 0.324 ;
        RECT 3.192 -0.048 3.288 0.216 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.048 0.684 4.392 0.756 ;
      RECT 4.32 0.108 4.392 0.756 ;
      RECT 4.32 0.396 4.7 0.468 ;
      RECT 4.048 0.108 4.392 0.18 ;
      RECT 2.88 0.108 2.952 0.72 ;
      RECT 2.88 0.508 3.6 0.58 ;
      RECT 3.528 0.396 3.6 0.58 ;
      RECT 3.312 0.396 3.384 0.58 ;
      RECT 3.528 0.396 4.032 0.468 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 3.096 0.108 3.168 0.364 ;
      RECT 3.096 0.108 3.492 0.18 ;
      RECT 2.008 0.656 2.592 0.728 ;
      RECT 2.52 0.252 2.592 0.728 ;
      RECT 2.008 0.5 2.08 0.728 ;
      RECT 2.34 0.252 2.592 0.324 ;
      RECT 2.34 0.156 2.412 0.324 ;
      RECT 2.16 0.512 2.324 0.584 ;
      RECT 2.16 0.328 2.232 0.584 ;
      RECT 2.088 0.108 2.16 0.4 ;
      RECT 1.584 0.108 2.16 0.18 ;
      RECT 1.8 0.252 1.872 0.628 ;
      RECT 1.74 0.348 1.964 0.42 ;
      RECT 1.74 0.252 1.888 0.42 ;
      RECT 1.228 0.684 1.548 0.756 ;
      RECT 1.228 0.108 1.3 0.756 ;
      RECT 1.112 0.108 1.3 0.18 ;
      RECT 0.484 0.396 0.792 0.468 ;
      RECT 0.72 0.108 0.792 0.468 ;
      RECT 0.18 0.108 0.792 0.18 ;
      RECT 2.664 0.376 2.736 0.58 ;
      RECT 1.58 0.368 1.652 0.552 ;
      RECT 1.372 0.232 1.444 0.54 ;
      RECT 0.864 0.332 0.936 0.488 ;
    LAYER M2 ;
      RECT 0.844 0.396 2.756 0.468 ;
      RECT 0.7 0.252 1.896 0.324 ;
      RECT 1.12 0.108 1.76 0.18 ;
    LAYER V1 ;
      RECT 2.664 0.396 2.736 0.468 ;
      RECT 1.804 0.252 1.876 0.324 ;
      RECT 1.668 0.108 1.74 0.18 ;
      RECT 1.58 0.396 1.652 0.468 ;
      RECT 1.372 0.252 1.444 0.324 ;
      RECT 1.12 0.108 1.192 0.18 ;
      RECT 0.864 0.396 0.936 0.468 ;
      RECT 0.72 0.252 0.792 0.324 ;
  END
END DFFLQx4_ASAP7_6t_fix

MACRO DHLx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.36 0.464 ;
        RECT 0.072 0.108 0.36 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.348 0.36 0.42 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.036 0.684 1.28 0.756 ;
        RECT 1.152 0.168 1.224 0.756 ;
      LAYER V0 ;
        RECT 1.152 0.392 1.224 0.464 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.684 3.168 0.756 ;
        RECT 3.096 0.108 3.168 0.756 ;
        RECT 2.988 0.108 3.168 0.18 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.88 0.252 2.952 0.488 ;
      RECT 2.84 0.252 2.952 0.324 ;
      RECT 2.3 0.684 2.74 0.756 ;
      RECT 2.66 0.108 2.74 0.756 ;
      RECT 2.016 0.108 2.088 0.36 ;
      RECT 2.016 0.108 2.74 0.18 ;
      RECT 2.412 0.54 2.56 0.612 ;
      RECT 2.412 0.376 2.484 0.612 ;
      RECT 1.476 0.684 1.86 0.756 ;
      RECT 1.788 0.108 1.86 0.756 ;
      RECT 1.788 0.516 2.304 0.588 ;
      RECT 2.232 0.28 2.304 0.588 ;
      RECT 1.508 0.108 1.86 0.18 ;
      RECT 1.584 0.252 1.656 0.46 ;
      RECT 1.508 0.252 1.656 0.324 ;
      RECT 1.368 0.54 1.56 0.612 ;
      RECT 1.368 0.392 1.44 0.612 ;
      RECT 0.592 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.592 0.108 0.936 0.18 ;
      RECT 0.592 0.54 0.792 0.612 ;
      RECT 0.72 0.324 0.792 0.612 ;
      RECT 0.552 0.324 0.792 0.396 ;
      RECT 0.088 0.54 0.212 0.612 ;
    LAYER M2 ;
      RECT 1.768 0.252 2.968 0.324 ;
      RECT 0.076 0.54 2.58 0.612 ;
      RECT 0.844 0.252 1.644 0.324 ;
    LAYER V1 ;
      RECT 2.872 0.252 2.944 0.324 ;
      RECT 2.472 0.54 2.544 0.612 ;
      RECT 1.788 0.252 1.86 0.324 ;
      RECT 1.552 0.252 1.624 0.324 ;
      RECT 1.376 0.54 1.448 0.612 ;
      RECT 0.864 0.252 0.936 0.324 ;
      RECT 0.612 0.54 0.684 0.612 ;
      RECT 0.096 0.54 0.168 0.612 ;
  END
END DHLx1_ASAP7_6t_fix

MACRO DHLx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx2_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.36 0.46 ;
        RECT 0.072 0.108 0.36 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.324 0.36 0.396 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.036 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 1.036 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.964 0.684 3.416 0.756 ;
        RECT 3.344 0.108 3.416 0.756 ;
        RECT 2.828 0.108 3.416 0.18 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.092 0.252 3.164 0.488 ;
      RECT 3.092 0.252 3.244 0.324 ;
      RECT 2.88 0.252 2.952 0.488 ;
      RECT 2.804 0.252 2.952 0.324 ;
      RECT 2.32 0.684 2.704 0.756 ;
      RECT 2.632 0.108 2.704 0.756 ;
      RECT 2.016 0.108 2.088 0.384 ;
      RECT 2.016 0.108 2.704 0.18 ;
      RECT 2.384 0.54 2.532 0.612 ;
      RECT 2.44 0.444 2.512 0.612 ;
      RECT 1.364 0.684 1.872 0.756 ;
      RECT 1.8 0.108 1.872 0.756 ;
      RECT 1.8 0.576 2.18 0.648 ;
      RECT 2.108 0.464 2.18 0.648 ;
      RECT 2.108 0.464 2.304 0.536 ;
      RECT 2.232 0.316 2.304 0.536 ;
      RECT 1.652 0.108 1.872 0.18 ;
      RECT 1.584 0.252 1.656 0.488 ;
      RECT 1.544 0.252 1.696 0.324 ;
      RECT 1.364 0.54 1.512 0.612 ;
      RECT 1.368 0.328 1.44 0.612 ;
      RECT 0.552 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.592 0.108 0.936 0.18 ;
      RECT 0.592 0.54 0.792 0.612 ;
      RECT 0.72 0.324 0.792 0.612 ;
      RECT 0.552 0.324 0.792 0.396 ;
      RECT 0.088 0.54 0.212 0.612 ;
    LAYER M2 ;
      RECT 1.78 0.252 3.192 0.324 ;
      RECT 0.076 0.54 2.532 0.612 ;
      RECT 0.844 0.252 1.648 0.324 ;
    LAYER V1 ;
      RECT 3.1 0.252 3.172 0.324 ;
      RECT 2.872 0.252 2.944 0.324 ;
      RECT 2.44 0.54 2.512 0.612 ;
      RECT 1.8 0.252 1.872 0.324 ;
      RECT 1.556 0.252 1.628 0.324 ;
      RECT 1.376 0.54 1.448 0.612 ;
      RECT 0.864 0.252 0.936 0.324 ;
      RECT 0.612 0.54 0.684 0.612 ;
      RECT 0.096 0.54 0.168 0.612 ;
  END
END DHLx2_ASAP7_6t_fix

MACRO DHLx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx3_ASAP7_6t_fix 0 0 ;
  SIZE 3.672 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.36 0.46 ;
        RECT 0.068 0.108 0.36 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.324 0.36 0.396 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.036 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 1.036 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.152 0.392 1.224 0.464 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.752 0.684 3.624 0.756 ;
        RECT 3.552 0.108 3.624 0.756 ;
        RECT 2.752 0.108 3.624 0.18 ;
      LAYER V0 ;
        RECT 2.772 0.684 2.844 0.756 ;
        RECT 2.772 0.108 2.844 0.18 ;
        RECT 3.204 0.684 3.276 0.756 ;
        RECT 3.204 0.108 3.276 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.672 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.672 0.912 ;
        RECT 3.408 0.54 3.504 0.912 ;
        RECT 2.976 0.54 3.072 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.672 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.672 0.048 ;
        RECT 3.408 -0.048 3.504 0.324 ;
        RECT 2.976 -0.048 3.072 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.304 0.252 3.376 0.484 ;
      RECT 3.304 0.252 3.452 0.324 ;
      RECT 3.088 0.252 3.16 0.484 ;
      RECT 3.012 0.252 3.16 0.324 ;
      RECT 2.832 0.252 2.904 0.484 ;
      RECT 2.756 0.252 2.904 0.324 ;
      RECT 2.3 0.684 2.644 0.756 ;
      RECT 2.572 0.108 2.644 0.756 ;
      RECT 2.016 0.108 2.088 0.404 ;
      RECT 2.016 0.108 2.644 0.18 ;
      RECT 2.352 0.54 2.5 0.612 ;
      RECT 2.428 0.392 2.5 0.612 ;
      RECT 1.364 0.684 1.872 0.756 ;
      RECT 1.8 0.108 1.872 0.756 ;
      RECT 1.652 0.108 1.872 0.18 ;
      RECT 1.584 0.252 1.656 0.492 ;
      RECT 1.508 0.252 1.656 0.324 ;
      RECT 1.364 0.54 1.512 0.612 ;
      RECT 1.368 0.38 1.44 0.612 ;
      RECT 0.592 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.592 0.108 0.936 0.18 ;
      RECT 0.592 0.54 0.792 0.612 ;
      RECT 0.72 0.324 0.792 0.612 ;
      RECT 0.552 0.324 0.792 0.396 ;
      RECT 2.232 0.292 2.304 0.476 ;
      RECT 0.068 0.54 0.216 0.612 ;
    LAYER M2 ;
      RECT 1.78 0.252 3.404 0.324 ;
      RECT 0.076 0.54 2.496 0.612 ;
      RECT 1.8 0.396 2.304 0.468 ;
      RECT 0.844 0.252 1.656 0.324 ;
    LAYER V1 ;
      RECT 3.312 0.252 3.384 0.324 ;
      RECT 3.048 0.252 3.12 0.324 ;
      RECT 2.804 0.252 2.876 0.324 ;
      RECT 2.392 0.54 2.464 0.612 ;
      RECT 2.232 0.396 2.304 0.468 ;
      RECT 1.8 0.252 1.872 0.324 ;
      RECT 1.8 0.396 1.872 0.468 ;
      RECT 1.564 0.252 1.636 0.324 ;
      RECT 1.372 0.54 1.444 0.612 ;
      RECT 0.864 0.252 0.936 0.324 ;
      RECT 0.612 0.54 0.684 0.612 ;
      RECT 0.096 0.54 0.168 0.612 ;
  END
END DHLx3_ASAP7_6t_fix

MACRO DLLx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx1_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.36 0.756 ;
        RECT 0.288 0.404 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.444 0.36 0.516 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.368 0.18 ;
        RECT 1.152 0.108 1.224 0.496 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.684 3.168 0.756 ;
        RECT 3.096 0.108 3.168 0.756 ;
        RECT 2.948 0.108 3.168 0.18 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.88 0.252 2.952 0.464 ;
      RECT 2.804 0.252 2.952 0.324 ;
      RECT 2.556 0.108 2.628 0.724 ;
      RECT 1.996 0.272 2.16 0.344 ;
      RECT 2.088 0.108 2.16 0.344 ;
      RECT 2.088 0.108 2.628 0.18 ;
      RECT 1.4 0.684 1.872 0.756 ;
      RECT 1.8 0.108 1.872 0.756 ;
      RECT 1.8 0.436 2.304 0.508 ;
      RECT 2.232 0.28 2.304 0.508 ;
      RECT 1.652 0.108 1.872 0.18 ;
      RECT 1.584 0.252 1.656 0.584 ;
      RECT 1.508 0.252 1.656 0.324 ;
      RECT 1.292 0.54 1.44 0.612 ;
      RECT 1.368 0.4 1.44 0.612 ;
      RECT 0.592 0.684 1.008 0.756 ;
      RECT 0.936 0.108 1.008 0.756 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.572 0.252 0.644 0.556 ;
      RECT 0.572 0.252 0.812 0.324 ;
      RECT 2.376 0.392 2.448 0.624 ;
      RECT 0.076 0.252 0.252 0.324 ;
    LAYER M2 ;
      RECT 1.8 0.252 2.972 0.324 ;
      RECT 0.916 0.54 2.448 0.612 ;
      RECT 0.076 0.252 1.656 0.324 ;
    LAYER V1 ;
      RECT 2.864 0.252 2.936 0.324 ;
      RECT 2.376 0.54 2.448 0.612 ;
      RECT 1.8 0.252 1.872 0.324 ;
      RECT 1.552 0.252 1.624 0.324 ;
      RECT 1.34 0.54 1.412 0.612 ;
      RECT 0.936 0.54 1.008 0.612 ;
      RECT 0.72 0.252 0.792 0.324 ;
      RECT 0.096 0.252 0.168 0.324 ;
  END
END DLLx1_ASAP7_6t_fix

MACRO DLLx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx2_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.36 0.46 ;
        RECT 0.068 0.108 0.36 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.324 0.36 0.396 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.112 1.368 0.184 ;
        RECT 1.152 0.112 1.224 0.488 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.772 0.684 3.388 0.756 ;
        RECT 3.316 0.108 3.388 0.756 ;
        RECT 2.752 0.108 3.388 0.18 ;
      LAYER V0 ;
        RECT 2.772 0.684 2.844 0.756 ;
        RECT 2.772 0.108 2.844 0.18 ;
        RECT 3.204 0.684 3.276 0.756 ;
        RECT 3.204 0.108 3.276 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 2.976 0.54 3.072 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 2.976 -0.048 3.072 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.956 0.54 3.168 0.612 ;
      RECT 3.096 0.36 3.168 0.612 ;
      RECT 2.576 0.108 2.648 0.72 ;
      RECT 2.016 0.108 2.088 0.36 ;
      RECT 2.016 0.108 2.648 0.18 ;
      RECT 1.456 0.684 1.872 0.756 ;
      RECT 1.8 0.108 1.872 0.756 ;
      RECT 1.8 0.548 2.304 0.62 ;
      RECT 2.232 0.288 2.304 0.62 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 1.516 0.54 1.664 0.612 ;
      RECT 1.592 0.376 1.664 0.612 ;
      RECT 0.592 0.684 1.008 0.756 ;
      RECT 0.936 0.108 1.008 0.756 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.572 0.54 0.792 0.612 ;
      RECT 0.72 0.324 0.792 0.612 ;
      RECT 0.552 0.324 0.792 0.396 ;
      RECT 2.404 0.38 2.476 0.528 ;
      RECT 1.344 0.316 1.416 0.488 ;
      RECT 0.076 0.54 0.256 0.612 ;
    LAYER M2 ;
      RECT 1.78 0.54 3.2 0.612 ;
      RECT 0.916 0.396 2.496 0.468 ;
      RECT 0.076 0.54 1.656 0.612 ;
    LAYER V1 ;
      RECT 3.04 0.54 3.112 0.612 ;
      RECT 2.404 0.396 2.476 0.468 ;
      RECT 1.8 0.54 1.872 0.612 ;
      RECT 1.564 0.54 1.636 0.612 ;
      RECT 1.344 0.396 1.416 0.468 ;
      RECT 0.936 0.396 1.008 0.468 ;
      RECT 0.624 0.54 0.696 0.612 ;
      RECT 0.096 0.54 0.168 0.612 ;
  END
END DLLx2_ASAP7_6t_fix

MACRO DLLx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLLx3_ASAP7_6t_fix 0 0 ;
  SIZE 3.672 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.36 0.46 ;
        RECT 0.068 0.108 0.36 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.324 0.36 0.396 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.444 0.18 ;
        RECT 1.152 0.108 1.224 0.552 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.684 3.604 0.756 ;
        RECT 3.528 0.144 3.604 0.756 ;
        RECT 2.968 0.144 3.604 0.216 ;
      LAYER V0 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.144 3.06 0.216 ;
        RECT 3.42 0.684 3.492 0.756 ;
        RECT 3.42 0.144 3.492 0.216 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.672 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.672 0.912 ;
        RECT 3.192 0.54 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.672 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.672 0.048 ;
        RECT 3.192 -0.048 3.288 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.112 -0.048 2.208 0.216 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.02 0.54 3.168 0.612 ;
      RECT 3.096 0.36 3.168 0.612 ;
      RECT 2.576 0.108 2.648 0.72 ;
      RECT 2.016 0.108 2.088 0.36 ;
      RECT 2.016 0.108 2.648 0.18 ;
      RECT 1.456 0.684 1.872 0.756 ;
      RECT 1.8 0.108 1.872 0.756 ;
      RECT 1.8 0.54 2.304 0.612 ;
      RECT 2.232 0.288 2.304 0.612 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 1.516 0.54 1.664 0.612 ;
      RECT 1.592 0.376 1.664 0.612 ;
      RECT 0.592 0.684 1.008 0.756 ;
      RECT 0.936 0.108 1.008 0.756 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.54 0.792 0.612 ;
      RECT 0.72 0.328 0.792 0.612 ;
      RECT 0.552 0.328 0.792 0.4 ;
      RECT 2.404 0.364 2.476 0.528 ;
      RECT 1.344 0.324 1.416 0.552 ;
      RECT 0.072 0.54 0.256 0.612 ;
    LAYER M2 ;
      RECT 1.8 0.54 3.2 0.612 ;
      RECT 0.916 0.396 2.496 0.468 ;
      RECT 0.076 0.54 1.656 0.612 ;
    LAYER V1 ;
      RECT 3.064 0.54 3.136 0.612 ;
      RECT 2.404 0.396 2.476 0.468 ;
      RECT 1.8 0.54 1.872 0.612 ;
      RECT 1.564 0.54 1.636 0.612 ;
      RECT 1.344 0.396 1.416 0.468 ;
      RECT 0.936 0.396 1.008 0.468 ;
      RECT 0.636 0.54 0.708 0.612 ;
      RECT 0.096 0.54 0.168 0.612 ;
  END
END DLLx3_ASAP7_6t_fix

MACRO FAx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAx1_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.144 0.38 2.304 0.452 ;
        RECT 2.144 0.26 2.216 0.452 ;
        RECT 1.588 0.26 2.216 0.332 ;
        RECT 1.864 0.108 2.012 0.332 ;
        RECT 0.72 0.54 1.66 0.612 ;
        RECT 1.588 0.26 1.66 0.612 ;
        RECT 0.788 0.684 1.008 0.756 ;
        RECT 0.936 0.54 1.008 0.756 ;
        RECT 0.72 0.396 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
        RECT 1.588 0.408 1.66 0.48 ;
        RECT 2.232 0.38 2.304 0.452 ;
    END
  END CI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.468 0.756 ;
        RECT 0.072 0.108 0.468 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 2.976 0.54 3.072 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 2.976 -0.048 3.072 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.296 0.54 1.988 0.612 ;
      LAYER M1 ;
        RECT 1.908 0.54 2.76 0.612 ;
        RECT 2.688 0.376 2.76 0.612 ;
        RECT 1.908 0.404 1.98 0.612 ;
        RECT 1.76 0.404 1.98 0.476 ;
        RECT 0.288 0.54 0.436 0.612 ;
        RECT 0.288 0.396 0.36 0.612 ;
      LAYER V1 ;
        RECT 0.296 0.54 0.368 0.612 ;
        RECT 1.916 0.54 1.988 0.612 ;
      LAYER V0 ;
        RECT 0.288 0.396 0.36 0.468 ;
        RECT 1.836 0.404 1.908 0.476 ;
        RECT 2.688 0.396 2.76 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.288 0.252 2.984 0.324 ;
      LAYER M1 ;
        RECT 2.98 0.252 3.052 0.48 ;
        RECT 2.904 0.252 3.052 0.324 ;
        RECT 1.324 0.396 1.488 0.468 ;
        RECT 1.324 0.252 1.396 0.468 ;
        RECT 0.94 0.252 1.396 0.324 ;
        RECT 0.94 0.108 1.012 0.324 ;
        RECT 0.592 0.108 1.012 0.18 ;
        RECT 0.504 0.252 0.664 0.324 ;
        RECT 0.592 0.108 0.664 0.324 ;
        RECT 0.504 0.252 0.576 0.42 ;
      LAYER V1 ;
        RECT 1.288 0.252 1.36 0.324 ;
        RECT 2.912 0.252 2.984 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.348 0.576 0.42 ;
        RECT 1.396 0.396 1.468 0.468 ;
        RECT 2.98 0.388 3.052 0.46 ;
    END
  END B
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.004 0.396 2.54 0.468 ;
      LAYER M1 ;
        RECT 2.428 0.396 2.576 0.468 ;
        RECT 0.936 0.396 1.084 0.468 ;
      LAYER V1 ;
        RECT 1.004 0.396 1.076 0.468 ;
        RECT 2.448 0.396 2.52 0.468 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
        RECT 2.448 0.396 2.52 0.468 ;
    END
  END CON
  OBS
    LAYER M1 ;
      RECT 2.092 0.684 3.332 0.756 ;
      RECT 2.124 0.108 3.276 0.18 ;
      RECT 1.24 0.684 1.784 0.756 ;
      RECT 1.26 0.108 1.764 0.18 ;
  END
END FAx1_ASAP7_6t_fix

MACRO FILLER_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER_ASAP7_6t_fix 0 0 ;
  SIZE 0.432 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.432 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.432 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.432 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.432 0.048 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
    END
  END VSS
END FILLER_ASAP7_6t_fix

MACRO FILLERxp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLERxp5_ASAP7_6t_fix 0 0 ;
  SIZE 0.216 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.216 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.216 0.912 ;
      LAYER V0 ;
        RECT 0.072 0.828 0.144 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.216 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.216 0.048 ;
      LAYER V0 ;
        RECT 0.072 -0.036 0.144 0.036 ;
    END
  END VSS
END FILLERxp5_ASAP7_6t_fix

MACRO HAx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HAx1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 1.344 0.756 ;
        RECT 0.472 0.252 0.544 0.756 ;
        RECT 0.396 0.252 0.544 0.324 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.252 0.468 0.324 ;
        RECT 1.044 0.684 1.116 0.756 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.328 0.648 2.424 0.912 ;
        RECT 1.896 0.648 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.692 0.396 2.116 0.468 ;
      LAYER M1 ;
        RECT 2.016 0.396 2.312 0.468 ;
        RECT 2.016 0.396 2.088 0.584 ;
        RECT 1.292 0.396 1.468 0.468 ;
        RECT 0.644 0.396 0.812 0.468 ;
      LAYER V1 ;
        RECT 0.712 0.396 0.784 0.468 ;
        RECT 1.3 0.396 1.372 0.468 ;
        RECT 2.024 0.396 2.096 0.468 ;
      LAYER V0 ;
        RECT 0.712 0.396 0.784 0.468 ;
        RECT 1.396 0.396 1.468 0.468 ;
        RECT 2.124 0.396 2.196 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.928 0.252 2.136 0.324 ;
      LAYER M1 ;
        RECT 1.872 0.252 2.312 0.324 ;
        RECT 1.872 0.252 1.944 0.576 ;
        RECT 1.8 0.412 1.944 0.484 ;
        RECT 0.956 0.396 1.104 0.468 ;
        RECT 0.956 0.252 1.028 0.468 ;
        RECT 0.88 0.252 1.028 0.324 ;
      LAYER V1 ;
        RECT 0.948 0.252 1.02 0.324 ;
        RECT 2.024 0.252 2.096 0.324 ;
      LAYER V0 ;
        RECT 1.032 0.396 1.104 0.468 ;
        RECT 1.8 0.412 1.872 0.484 ;
    END
  END B
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.196 0.54 1.684 0.612 ;
      LAYER M1 ;
        RECT 1.584 0.684 2.304 0.756 ;
        RECT 1.58 0.252 1.748 0.324 ;
        RECT 1.584 0.252 1.656 0.756 ;
        RECT 0.216 0.396 0.288 0.728 ;
        RECT 0.072 0.396 0.288 0.468 ;
      LAYER V1 ;
        RECT 0.216 0.54 0.288 0.612 ;
        RECT 1.584 0.54 1.656 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 1.656 0.252 1.728 0.324 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 2.124 0.684 2.196 0.756 ;
    END
  END CON
  OBS
    LAYER M1 ;
      RECT 2.124 0.108 2.412 0.18 ;
      RECT 1.476 0.108 2 0.18 ;
      RECT 0.656 0.54 1.368 0.612 ;
      RECT 0.16 0.108 1.332 0.18 ;
    LAYER M2 ;
      RECT 1.232 0.108 2.412 0.18 ;
    LAYER V1 ;
      RECT 2.252 0.108 2.324 0.18 ;
      RECT 1.252 0.108 1.324 0.18 ;
  END
END HAx1_ASAP7_6t_fix

MACRO HAxp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HAxp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.348 0.396 1.572 0.468 ;
        RECT 1.5 0.252 1.572 0.468 ;
        RECT 0.848 0.252 1.572 0.324 ;
        RECT 0.848 0.108 0.92 0.324 ;
        RECT 0.072 0.108 0.92 0.18 ;
        RECT 0.072 0.684 0.224 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.576 0.396 1.148 0.468 ;
        RECT 0.576 0.54 0.812 0.612 ;
        RECT 0.576 0.396 0.648 0.612 ;
      LAYER V0 ;
        RECT 1.04 0.396 1.112 0.468 ;
    END
  END B
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.724 0.612 ;
        RECT 1.652 0.38 1.724 0.612 ;
        RECT 0.36 0.684 1.008 0.756 ;
        RECT 0.936 0.54 1.008 0.756 ;
        RECT 0.36 0.252 0.508 0.324 ;
        RECT 0.36 0.252 0.432 0.756 ;
      LAYER V0 ;
        RECT 0.36 0.524 0.432 0.596 ;
        RECT 0.436 0.252 0.508 0.324 ;
        RECT 1.652 0.4 1.724 0.472 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.692 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.044 0.108 1.548 0.18 ;
  END
END HAxp5_ASAP7_6t_fix

MACRO HB1xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB1xp67_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.208 0.684 0.36 0.756 ;
        RECT 0.288 0.108 0.36 0.756 ;
        RECT 0.208 0.108 0.36 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.284 0.36 0.356 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.684 0.792 0.756 ;
        RECT 0.72 0.108 0.792 0.756 ;
        RECT 0.612 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
END HB1xp67_ASAP7_6t_fix

MACRO HB2xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB2xp67_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.6 -0.048 0.696 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.808 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.576 0.756 ;
      RECT 0.504 0.108 0.576 0.756 ;
      RECT 0.504 0.392 0.812 0.464 ;
      RECT 0.396 0.108 0.576 0.18 ;
  END
END HB2xp67_ASAP7_6t_fix

MACRO HB3xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB3xp67_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.388 0.416 0.46 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.388 0.36 0.46 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 1.024 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.684 0.792 0.756 ;
      RECT 0.72 0.108 0.792 0.756 ;
      RECT 0.72 0.388 1.028 0.46 ;
      RECT 0.612 0.108 0.792 0.18 ;
  END
END HB3xp67_ASAP7_6t_fix

MACRO HB4xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB4xp67_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.388 0.444 0.46 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.288 0.388 0.36 0.46 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 1.24 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.684 0.792 0.756 ;
      RECT 0.72 0.108 0.792 0.756 ;
      RECT 0.72 0.388 1.244 0.46 ;
      RECT 0.612 0.108 0.792 0.18 ;
  END
END HB4xp67_ASAP7_6t_fix

MACRO ICGx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx1_ASAP7_6t_fix 0 0 ;
  SIZE 4.104 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.308 0.468 ;
        RECT 0.072 0.108 0.232 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.216 0.396 0.288 0.468 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 3.74 0.684 4.032 0.756 ;
        RECT 3.96 0.108 4.032 0.756 ;
        RECT 3.74 0.108 4.032 0.18 ;
      LAYER V0 ;
        RECT 3.852 0.684 3.924 0.756 ;
        RECT 3.852 0.108 3.924 0.18 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.54 0.576 0.612 ;
        RECT 0.504 0.28 0.576 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.104 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.104 0.912 ;
        RECT 3.624 0.54 3.72 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 1.896 0.648 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.104 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.104 0.048 ;
        RECT 3.624 -0.048 3.72 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 1.896 -0.048 1.992 0.216 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
    END
  END VSS
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 2.66 0.54 3.292 0.612 ;
        RECT 0.916 0.396 2.688 0.468 ;
      LAYER M1 ;
        RECT 3.2 0.472 3.272 0.62 ;
        RECT 2.52 0.54 2.76 0.612 ;
        RECT 2.52 0.396 2.74 0.468 ;
        RECT 2.52 0.396 2.592 0.612 ;
        RECT 1.584 0.28 1.656 0.584 ;
        RECT 0.936 0.136 1.008 0.48 ;
      LAYER V1 ;
        RECT 0.936 0.396 1.008 0.468 ;
        RECT 1.584 0.396 1.656 0.468 ;
        RECT 2.528 0.396 2.6 0.468 ;
        RECT 2.68 0.54 2.752 0.612 ;
        RECT 3.2 0.54 3.272 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.388 1.008 0.46 ;
        RECT 1.584 0.396 1.656 0.468 ;
        RECT 2.648 0.396 2.72 0.468 ;
        RECT 3.2 0.496 3.272 0.568 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 3.4 0.684 3.6 0.756 ;
      RECT 3.528 0.54 3.6 0.756 ;
      RECT 3.528 0.54 3.816 0.612 ;
      RECT 3.744 0.252 3.816 0.612 ;
      RECT 3.184 0.252 3.816 0.324 ;
      RECT 1.012 0.684 1.872 0.756 ;
      RECT 1.8 0.512 1.872 0.756 ;
      RECT 1.296 0.108 1.368 0.756 ;
      RECT 1.8 0.512 2.108 0.584 ;
      RECT 2.88 0.108 2.952 0.48 ;
      RECT 1.296 0.108 2.952 0.18 ;
      RECT 2.376 0.684 2.66 0.756 ;
      RECT 2.376 0.252 2.448 0.756 ;
      RECT 2.376 0.252 2.636 0.324 ;
      RECT 2.04 0.684 2.304 0.756 ;
      RECT 2.228 0.28 2.304 0.756 ;
      RECT 1.78 0.28 2.304 0.352 ;
      RECT 1.076 0.54 1.224 0.612 ;
      RECT 1.152 0.324 1.224 0.612 ;
      RECT 0.148 0.684 0.792 0.756 ;
      RECT 0.72 0.108 0.792 0.756 ;
      RECT 0.356 0.108 0.792 0.18 ;
      RECT 3.444 0.396 3.596 0.468 ;
      RECT 2.932 0.684 3.08 0.756 ;
    LAYER M2 ;
      RECT 2.86 0.396 3.604 0.468 ;
      RECT 2.956 0.684 3.5 0.756 ;
      RECT 1.124 0.54 2.468 0.612 ;
    LAYER V1 ;
      RECT 3.512 0.396 3.584 0.468 ;
      RECT 3.408 0.684 3.48 0.756 ;
      RECT 2.976 0.684 3.048 0.756 ;
      RECT 2.88 0.396 2.952 0.468 ;
      RECT 2.376 0.54 2.448 0.612 ;
      RECT 1.144 0.54 1.216 0.612 ;
  END
END ICGx1_ASAP7_6t_fix

MACRO ICGx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx2_ASAP7_6t_fix 0 0 ;
  SIZE 4.32 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.308 0.468 ;
        RECT 0.072 0.108 0.232 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.216 0.396 0.288 0.468 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 3.74 0.684 4.248 0.756 ;
        RECT 4.176 0.108 4.248 0.756 ;
        RECT 3.74 0.108 4.248 0.18 ;
      LAYER V0 ;
        RECT 3.852 0.684 3.924 0.756 ;
        RECT 3.852 0.108 3.924 0.18 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.54 0.576 0.612 ;
        RECT 0.504 0.28 0.576 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.32 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.32 0.912 ;
        RECT 4.056 0.54 4.152 0.912 ;
        RECT 3.624 0.54 3.72 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 1.896 0.648 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.32 0.048 ;
        RECT 4.056 -0.048 4.152 0.324 ;
        RECT 3.624 -0.048 3.72 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 1.896 -0.048 1.992 0.216 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
    END
  END VSS
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 2.66 0.54 3.292 0.612 ;
        RECT 0.916 0.396 2.688 0.468 ;
      LAYER M1 ;
        RECT 3.2 0.472 3.272 0.62 ;
        RECT 2.52 0.54 2.76 0.612 ;
        RECT 2.52 0.396 2.74 0.468 ;
        RECT 2.52 0.396 2.592 0.612 ;
        RECT 1.584 0.28 1.656 0.584 ;
        RECT 0.936 0.136 1.008 0.48 ;
      LAYER V1 ;
        RECT 0.936 0.396 1.008 0.468 ;
        RECT 1.584 0.396 1.656 0.468 ;
        RECT 2.528 0.396 2.6 0.468 ;
        RECT 2.68 0.54 2.752 0.612 ;
        RECT 3.2 0.54 3.272 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.388 1.008 0.46 ;
        RECT 1.584 0.396 1.656 0.468 ;
        RECT 2.648 0.396 2.72 0.468 ;
        RECT 3.2 0.496 3.272 0.568 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 3.4 0.684 3.6 0.756 ;
      RECT 3.528 0.54 3.6 0.756 ;
      RECT 3.528 0.54 3.816 0.612 ;
      RECT 3.744 0.252 3.816 0.612 ;
      RECT 3.184 0.252 3.816 0.324 ;
      RECT 1.012 0.684 1.872 0.756 ;
      RECT 1.8 0.512 1.872 0.756 ;
      RECT 1.296 0.108 1.368 0.756 ;
      RECT 1.8 0.512 2.108 0.584 ;
      RECT 2.88 0.108 2.952 0.48 ;
      RECT 1.296 0.108 2.952 0.18 ;
      RECT 2.376 0.684 2.66 0.756 ;
      RECT 2.376 0.252 2.448 0.756 ;
      RECT 2.376 0.252 2.636 0.324 ;
      RECT 2.04 0.684 2.304 0.756 ;
      RECT 2.228 0.28 2.304 0.756 ;
      RECT 1.78 0.28 2.304 0.352 ;
      RECT 1.076 0.54 1.224 0.612 ;
      RECT 1.152 0.324 1.224 0.612 ;
      RECT 0.148 0.684 0.792 0.756 ;
      RECT 0.72 0.108 0.792 0.756 ;
      RECT 0.356 0.108 0.792 0.18 ;
      RECT 3.444 0.396 3.596 0.468 ;
      RECT 2.932 0.684 3.08 0.756 ;
    LAYER M2 ;
      RECT 2.86 0.396 3.604 0.468 ;
      RECT 2.956 0.684 3.5 0.756 ;
      RECT 1.124 0.54 2.468 0.612 ;
    LAYER V1 ;
      RECT 3.512 0.396 3.584 0.468 ;
      RECT 3.408 0.684 3.48 0.756 ;
      RECT 2.976 0.684 3.048 0.756 ;
      RECT 2.88 0.396 2.952 0.468 ;
      RECT 2.376 0.54 2.448 0.612 ;
      RECT 1.144 0.54 1.216 0.612 ;
  END
END ICGx2_ASAP7_6t_fix

MACRO ICGx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGx3_ASAP7_6t_fix 0 0 ;
  SIZE 4.536 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.308 0.468 ;
        RECT 0.072 0.108 0.232 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.216 0.396 0.288 0.468 ;
    END
  END ENA
  PIN GCLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 3.74 0.684 4.464 0.756 ;
        RECT 4.392 0.108 4.464 0.756 ;
        RECT 3.74 0.108 4.464 0.18 ;
      LAYER V0 ;
        RECT 3.852 0.684 3.924 0.756 ;
        RECT 3.852 0.108 3.924 0.18 ;
        RECT 4.284 0.684 4.356 0.756 ;
        RECT 4.284 0.108 4.356 0.18 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.54 0.576 0.612 ;
        RECT 0.504 0.28 0.576 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.536 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.536 0.912 ;
        RECT 4.056 0.54 4.152 0.912 ;
        RECT 3.624 0.54 3.72 0.912 ;
        RECT 3.192 0.648 3.288 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 1.896 0.648 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.536 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.536 0.048 ;
        RECT 4.056 -0.048 4.152 0.324 ;
        RECT 3.624 -0.048 3.72 0.324 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 1.896 -0.048 1.992 0.216 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
    END
  END VSS
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 2.66 0.54 3.292 0.612 ;
        RECT 0.916 0.396 2.688 0.468 ;
      LAYER M1 ;
        RECT 3.2 0.472 3.272 0.62 ;
        RECT 2.52 0.54 2.76 0.612 ;
        RECT 2.52 0.396 2.74 0.468 ;
        RECT 2.52 0.396 2.592 0.612 ;
        RECT 1.584 0.28 1.656 0.584 ;
        RECT 0.936 0.136 1.008 0.48 ;
      LAYER V1 ;
        RECT 0.936 0.396 1.008 0.468 ;
        RECT 1.584 0.396 1.656 0.468 ;
        RECT 2.528 0.396 2.6 0.468 ;
        RECT 2.68 0.54 2.752 0.612 ;
        RECT 3.2 0.54 3.272 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.388 1.008 0.46 ;
        RECT 1.584 0.396 1.656 0.468 ;
        RECT 2.648 0.396 2.72 0.468 ;
        RECT 3.2 0.496 3.272 0.568 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 3.4 0.684 3.6 0.756 ;
      RECT 3.528 0.54 3.6 0.756 ;
      RECT 3.528 0.54 3.816 0.612 ;
      RECT 3.744 0.252 3.816 0.612 ;
      RECT 3.184 0.252 3.816 0.324 ;
      RECT 1.012 0.684 1.872 0.756 ;
      RECT 1.8 0.512 1.872 0.756 ;
      RECT 1.296 0.108 1.368 0.756 ;
      RECT 1.8 0.512 2.108 0.584 ;
      RECT 2.88 0.108 2.952 0.48 ;
      RECT 1.296 0.108 2.952 0.18 ;
      RECT 2.376 0.684 2.66 0.756 ;
      RECT 2.376 0.252 2.448 0.756 ;
      RECT 2.376 0.252 2.636 0.324 ;
      RECT 2.04 0.684 2.304 0.756 ;
      RECT 2.228 0.28 2.304 0.756 ;
      RECT 1.78 0.28 2.304 0.352 ;
      RECT 1.076 0.54 1.224 0.612 ;
      RECT 1.152 0.324 1.224 0.612 ;
      RECT 0.148 0.684 0.792 0.756 ;
      RECT 0.72 0.108 0.792 0.756 ;
      RECT 0.356 0.108 0.792 0.18 ;
      RECT 3.444 0.396 3.596 0.468 ;
      RECT 2.932 0.684 3.08 0.756 ;
    LAYER M2 ;
      RECT 2.86 0.396 3.604 0.468 ;
      RECT 2.956 0.684 3.5 0.756 ;
      RECT 1.124 0.54 2.468 0.612 ;
    LAYER V1 ;
      RECT 3.512 0.396 3.584 0.468 ;
      RECT 3.408 0.684 3.48 0.756 ;
      RECT 2.976 0.684 3.048 0.756 ;
      RECT 2.88 0.396 2.952 0.468 ;
      RECT 2.376 0.54 2.448 0.612 ;
      RECT 1.144 0.54 1.216 0.612 ;
  END
END ICGx3_ASAP7_6t_fix

MACRO INVx11_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx11_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 2.628 0.756 ;
        RECT 0.396 0.108 2.628 0.18 ;
        RECT 1.152 0.108 1.224 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
    END
  END Y
END INVx11_ASAP7_6t_fix

MACRO INVx13_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx13_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 3.06 0.756 ;
        RECT 0.396 0.108 3.06 0.18 ;
        RECT 1.152 0.108 1.224 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.988 0.684 3.06 0.756 ;
        RECT 2.988 0.108 3.06 0.18 ;
    END
  END Y
END INVx13_ASAP7_6t_fix

MACRO INVx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1_ASAP7_6t_fix 0 0 ;
  SIZE 0.648 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.648 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.648 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.648 0.048 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 0.584 0.756 ;
        RECT 0.396 0.108 0.584 0.18 ;
        RECT 0.504 0.108 0.576 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
END INVx1_ASAP7_6t_fix

MACRO INVx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 0.728 0.756 ;
        RECT 0.396 0.108 0.728 0.18 ;
        RECT 0.648 0.108 0.72 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
END INVx2_ASAP7_6t_fix

MACRO INVx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx3_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 0.9 0.756 ;
        RECT 0.396 0.108 0.9 0.18 ;
        RECT 0.504 0.108 0.576 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
END INVx3_ASAP7_6t_fix

MACRO INVx4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.396 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
END INVx4_ASAP7_6t_fix

MACRO INVx5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx5_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 1.368 0.756 ;
        RECT 0.396 0.108 1.368 0.18 ;
        RECT 1.152 0.108 1.224 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
END INVx5_ASAP7_6t_fix

MACRO INVx6_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx6_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 1.332 0.756 ;
        RECT 0.396 0.108 1.332 0.18 ;
        RECT 1.044 0.108 1.116 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
    END
  END Y
END INVx6_ASAP7_6t_fix

MACRO INVx8_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.22 0.756 ;
        RECT 0.064 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 1.764 0.756 ;
        RECT 0.396 0.108 1.764 0.18 ;
        RECT 1.152 0.108 1.224 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
END INVx8_ASAP7_6t_fix

MACRO INVxp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp33_ASAP7_6t_fix 0 0 ;
  SIZE 0.648 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.648 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.648 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.648 0.048 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 0.576 0.756 ;
        RECT 0.504 0.108 0.576 0.756 ;
        RECT 0.396 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
END INVxp33_ASAP7_6t_fix

MACRO INVxp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVxp67_ASAP7_6t_fix 0 0 ;
  SIZE 0.648 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.36 0.612 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.648 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.648 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.648 0.048 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.684 0.576 0.756 ;
        RECT 0.504 0.108 0.576 0.756 ;
        RECT 0.396 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
END INVxp67_ASAP7_6t_fix

MACRO MAJIxp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJIxp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.54 1.444 0.612 ;
        RECT 1.296 0.252 1.444 0.324 ;
        RECT 1.296 0.252 1.368 0.612 ;
      LAYER V0 ;
        RECT 1.296 0.396 1.368 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.712 0.396 0.98 0.468 ;
        RECT 0.072 0.54 0.784 0.612 ;
        RECT 0.712 0.392 0.784 0.612 ;
        RECT 0.072 0.396 0.332 0.468 ;
        RECT 0.072 0.396 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.24 0.396 0.312 0.468 ;
        RECT 0.908 0.396 0.98 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.456 0.384 0.604 0.456 ;
        RECT 0.456 0.252 0.528 0.456 ;
        RECT 0.192 0.252 0.528 0.324 ;
        RECT 0.192 0.108 0.264 0.324 ;
        RECT 0.064 0.108 0.264 0.18 ;
      LAYER V0 ;
        RECT 0.532 0.384 0.604 0.456 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.54 1.152 0.612 ;
        RECT 1.08 0.252 1.152 0.612 ;
        RECT 0.908 0.252 1.152 0.324 ;
      LAYER V0 ;
        RECT 0.908 0.54 0.98 0.612 ;
        RECT 0.908 0.252 0.98 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 1.376 0.756 ;
      RECT 0.396 0.108 1.352 0.18 ;
  END
END MAJIxp5_ASAP7_6t_fix

MACRO MAJx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx2_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.228 0.612 ;
        RECT 0.072 0.252 0.228 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 1.388 0.756 ;
        RECT 1.24 0.54 1.312 0.756 ;
        RECT 0.936 0.54 1.312 0.612 ;
        RECT 0.936 0.396 1.008 0.612 ;
        RECT 0.852 0.396 1.008 0.468 ;
      LAYER V0 ;
        RECT 0.852 0.396 0.924 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.44 0.108 1.872 0.18 ;
        RECT 1.512 0.592 1.584 0.756 ;
      LAYER V0 ;
        RECT 1.476 0.108 1.548 0.18 ;
        RECT 1.512 0.612 1.584 0.684 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.508 0.396 1.272 0.468 ;
      LAYER M1 ;
        RECT 1.132 0.396 1.28 0.468 ;
        RECT 0.508 0.396 0.728 0.468 ;
      LAYER V1 ;
        RECT 0.532 0.396 0.604 0.468 ;
        RECT 1.152 0.396 1.224 0.468 ;
      LAYER V0 ;
        RECT 0.532 0.396 0.604 0.468 ;
        RECT 1.18 0.396 1.252 0.468 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.328 0.54 0.652 0.612 ;
      RECT 0.328 0.252 0.4 0.612 ;
      RECT 1.584 0.252 1.656 0.46 ;
      RECT 0.328 0.252 1.656 0.324 ;
      RECT 0.16 0.108 1.136 0.18 ;
      RECT 0.18 0.684 1.116 0.756 ;
  END
END MAJx2_ASAP7_6t_fix

MACRO MAJx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJx3_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.508 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.68 0.54 1.372 0.612 ;
        RECT 1.3 0.396 1.372 0.612 ;
        RECT 1.152 0.396 1.372 0.468 ;
        RECT 0.68 0.396 0.752 0.612 ;
        RECT 0.496 0.396 0.752 0.468 ;
      LAYER V0 ;
        RECT 0.528 0.396 0.6 0.468 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.884 0.396 1.66 0.468 ;
      LAYER M1 ;
        RECT 0.88 0.396 1.028 0.468 ;
      LAYER V1 ;
        RECT 0.908 0.396 0.98 0.468 ;
      LAYER V0 ;
        RECT 0.908 0.396 0.98 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.684 2.016 0.756 ;
        RECT 1.456 0.108 2.016 0.18 ;
        RECT 1.8 0.108 1.872 0.756 ;
      LAYER V0 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
        RECT 1.908 0.684 1.98 0.756 ;
        RECT 1.908 0.108 1.98 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.324 0.54 0.556 0.612 ;
      RECT 1.472 0.252 1.544 0.584 ;
      RECT 0.324 0.252 0.396 0.612 ;
      RECT 0.324 0.252 1.544 0.324 ;
      RECT 0.16 0.108 1.136 0.18 ;
      RECT 0.16 0.684 1.136 0.756 ;
  END
END MAJx3_ASAP7_6t_fix

MACRO MUX2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.684 2.38 0.756 ;
        RECT 2.232 0.252 2.38 0.324 ;
        RECT 2.232 0.252 2.304 0.756 ;
      LAYER V0 ;
        RECT 2.232 0.388 2.304 0.46 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.54 2.088 0.612 ;
        RECT 2.016 0.252 2.088 0.612 ;
        RECT 1.94 0.252 2.088 0.324 ;
      LAYER V0 ;
        RECT 2.016 0.388 2.088 0.46 ;
    END
  END B
  PIN O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.292 0.756 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.18 0.108 0.252 0.18 ;
    END
  END O
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 1.696 0.468 ;
        RECT 1.624 0.252 1.696 0.468 ;
        RECT 1.476 0.252 1.696 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
        RECT 1.44 0.396 1.512 0.468 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.564 0.54 1.84 0.612 ;
      RECT 1.768 0.108 1.84 0.612 ;
      RECT 1.044 0.108 2.412 0.18 ;
      RECT 0.288 0.54 1.332 0.612 ;
      RECT 0.288 0.252 0.36 0.612 ;
      RECT 0.288 0.252 1.332 0.324 ;
      RECT 1.044 0.684 1.98 0.756 ;
  END
END MUX2x1_ASAP7_6t_fix

MACRO MUX2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.396 1.452 0.468 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.54 1.948 0.612 ;
        RECT 1.8 0.252 1.872 0.612 ;
        RECT 1.712 0.252 1.872 0.324 ;
      LAYER V0 ;
        RECT 1.8 0.388 1.872 0.46 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.704 0.18 ;
        RECT 0.072 0.54 0.636 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.564 0.54 0.636 0.612 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.36 0.252 2.108 0.324 ;
      LAYER M1 ;
        RECT 2.36 0.396 2.592 0.468 ;
        RECT 2.52 0.252 2.592 0.468 ;
        RECT 2.028 0.252 2.592 0.324 ;
        RECT 0.372 0.252 0.52 0.324 ;
        RECT 0.296 0.396 0.444 0.468 ;
        RECT 0.372 0.252 0.444 0.468 ;
      LAYER V1 ;
        RECT 0.38 0.252 0.452 0.324 ;
        RECT 2.036 0.252 2.108 0.324 ;
      LAYER V0 ;
        RECT 0.296 0.396 0.368 0.468 ;
        RECT 2.448 0.396 2.52 0.468 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2.304 0.54 2.736 0.612 ;
      RECT 2.664 0.108 2.736 0.612 ;
      RECT 0.792 0.252 0.864 0.468 ;
      RECT 0.792 0.252 1.332 0.324 ;
      RECT 1.26 0.108 1.332 0.324 ;
      RECT 1.26 0.108 2.736 0.18 ;
      RECT 0.18 0.684 1.136 0.756 ;
      RECT 1.064 0.54 1.136 0.756 ;
      RECT 1.064 0.54 1.656 0.612 ;
      RECT 1.584 0.404 1.656 0.612 ;
      RECT 1.26 0.684 2.628 0.756 ;
      RECT 0.828 0.108 1.116 0.18 ;
  END
END MUX2x2_ASAP7_6t_fix

MACRO NAND2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.36 0.324 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.684 1.228 0.756 ;
        RECT 1.008 0.252 1.228 0.324 ;
        RECT 1.008 0.252 1.08 0.756 ;
        RECT 0.828 0.412 1.08 0.484 ;
      LAYER V0 ;
        RECT 0.828 0.412 0.9 0.484 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 0.9 0.756 ;
        RECT 0.576 0.252 0.9 0.324 ;
        RECT 0.576 0.252 0.648 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.252 0.9 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END NAND2x1_ASAP7_6t_fix

MACRO NAND2x1p5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1p5_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 1.136 0.468 ;
        RECT 0.428 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.044 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.252 1.332 0.324 ;
      RECT 0.396 0.108 0.9 0.18 ;
  END
END NAND2x1p5_ASAP7_6t_fix

MACRO NAND2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.252 1.24 0.324 ;
        RECT 0.856 0.396 1.08 0.468 ;
        RECT 1.008 0.252 1.08 0.468 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.464 0.396 1.764 0.468 ;
        RECT 0.62 0.54 1.536 0.612 ;
        RECT 1.464 0.396 1.536 0.612 ;
        RECT 0.62 0.396 0.692 0.612 ;
        RECT 0.216 0.396 0.692 0.468 ;
        RECT 0.064 0.684 0.288 0.756 ;
        RECT 0.216 0.396 0.288 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.396 0.468 0.468 ;
        RECT 1.692 0.396 1.764 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 2.088 0.756 ;
        RECT 2.016 0.252 2.088 0.756 ;
        RECT 1.692 0.252 2.088 0.324 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.252 1.764 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.252 0.144 0.496 ;
      RECT 0.072 0.252 0.468 0.324 ;
      RECT 0.16 0.108 2 0.18 ;
  END
END NAND2x2_ASAP7_6t_fix

MACRO NAND2xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp33_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.448 0.18 ;
        RECT 0.072 0.684 0.252 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.356 0.524 0.576 0.596 ;
        RECT 0.504 0.252 0.576 0.596 ;
        RECT 0.244 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.684 0.792 0.756 ;
        RECT 0.72 0.108 0.792 0.756 ;
        RECT 0.572 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.72 0.256 0.792 0.328 ;
    END
  END Y
END NAND2xp33_ASAP7_6t_fix

MACRO NAND2xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp5_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.368 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.368 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.684 0.792 0.756 ;
        RECT 0.72 0.108 0.792 0.756 ;
        RECT 0.612 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
END NAND2xp5_ASAP7_6t_fix

MACRO NAND2xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2xp67_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.224 0.756 ;
        RECT 0.072 0.252 0.224 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 0.936 0.468 ;
        RECT 0.424 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.424 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.396 0.9 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.684 1.224 0.756 ;
        RECT 1.152 0.252 1.224 0.756 ;
        RECT 0.828 0.252 1.224 0.324 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.828 0.252 0.9 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.108 1.116 0.18 ;
  END
END NAND2xp67_ASAP7_6t_fix

MACRO NAND3x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.684 2.304 0.756 ;
        RECT 2.016 0.396 2.304 0.468 ;
        RECT 2.016 0.396 2.088 0.756 ;
      LAYER V0 ;
        RECT 2.124 0.396 2.196 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 1.116 0.468 ;
        RECT 0.428 0.684 0.576 0.756 ;
        RECT 0.504 0.396 0.576 0.756 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
        RECT 0.16 0.108 0.704 0.18 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 0.168 -0.048 0.264 0.324 ;
        RECT 0.6 0.108 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.252 2.216 0.324 ;
        RECT 0.808 0.684 1.872 0.756 ;
        RECT 1.8 0.252 1.872 0.756 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.252 1.764 0.324 ;
        RECT 2.124 0.252 2.196 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.108 1.98 0.18 ;
      RECT 0.396 0.252 1.352 0.324 ;
  END
END NAND3x1_ASAP7_6t_fix

MACRO NAND3x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2_ASAP7_6t_fix 0 0 ;
  SIZE 4.32 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.904 0.396 3.148 0.468 ;
        RECT 1.132 0.54 2.976 0.612 ;
        RECT 2.904 0.396 2.976 0.612 ;
        RECT 1.132 0.396 1.204 0.612 ;
        RECT 0.828 0.396 1.204 0.468 ;
        RECT 0.828 0.28 0.9 0.468 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
        RECT 2.988 0.396 3.06 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.788 0.396 2.532 0.468 ;
      LAYER V0 ;
        RECT 2.124 0.396 2.196 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.32 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 4.32 0.912 ;
        RECT 3.408 0.54 3.504 0.912 ;
        RECT 2.976 0.54 3.072 0.912 ;
        RECT 2.544 0.54 2.64 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
        RECT 1.672 0.108 2.648 0.18 ;
      LAYER LISD ;
        RECT 0 -0.048 4.32 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 2.544 0.108 2.64 0.324 ;
        RECT 1.68 0.108 1.776 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.108 0.684 4.248 0.756 ;
        RECT 4.176 0.252 4.248 0.756 ;
        RECT 3.616 0.252 4.248 0.324 ;
        RECT 0.108 0.252 0.704 0.324 ;
        RECT 0.108 0.252 0.18 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.252 0.252 0.324 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.252 0.684 0.324 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 2.772 0.684 2.844 0.756 ;
        RECT 3.636 0.684 3.708 0.756 ;
        RECT 3.636 0.252 3.708 0.324 ;
        RECT 4.068 0.252 4.14 0.324 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.428 0.54 3.896 0.612 ;
      LAYER M1 ;
        RECT 3.724 0.54 3.888 0.612 ;
        RECT 3.724 0.396 3.796 0.612 ;
        RECT 3.552 0.396 3.796 0.468 ;
        RECT 0.284 0.54 0.6 0.612 ;
        RECT 0.284 0.396 0.6 0.468 ;
        RECT 0.284 0.396 0.356 0.612 ;
      LAYER V1 ;
        RECT 0.456 0.54 0.528 0.612 ;
        RECT 3.796 0.54 3.868 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.396 0.468 0.468 ;
        RECT 3.636 0.396 3.708 0.468 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 2.968 0.108 3.944 0.18 ;
      RECT 1.024 0.252 3.296 0.324 ;
      RECT 0.376 0.108 1.352 0.18 ;
  END
END NAND3x2_ASAP7_6t_fix

MACRO NAND3xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.108 0.552 0.18 ;
        RECT 0.256 0.54 0.404 0.612 ;
        RECT 0.288 0.108 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.288 0.396 0.36 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.54 0.792 0.612 ;
        RECT 0.504 0.252 0.792 0.324 ;
        RECT 0.504 0.252 0.576 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.676 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.684 0.756 ;
        RECT 0.072 0.28 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.612 0.684 0.684 0.756 ;
    END
  END Y
END NAND3xp33_ASAP7_6t_fix

MACRO NAND4xp25_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp25_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.54 1.224 0.612 ;
        RECT 1.008 0.108 1.224 0.18 ;
        RECT 1.008 0.108 1.08 0.612 ;
      LAYER V0 ;
        RECT 1.008 0.396 1.08 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 0.54 0.792 0.612 ;
        RECT 0.72 0.108 0.792 0.612 ;
        RECT 0.644 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.244 0.396 0.648 0.468 ;
        RECT 0.576 0.252 0.648 0.468 ;
        RECT 0.428 0.252 0.648 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.52 0.18 ;
        RECT 0.072 0.54 0.224 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.684 1.116 0.756 ;
        RECT 0.864 0.244 0.936 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 1.044 0.684 1.116 0.756 ;
    END
  END Y
END NAND4xp25_ASAP7_6t_fix

MACRO NAND4xp75_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4xp75_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.54 0.54 2.744 0.612 ;
        RECT 2.54 0.396 2.612 0.612 ;
        RECT 2.232 0.396 2.612 0.468 ;
      LAYER V0 ;
        RECT 2.34 0.396 2.412 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.396 2.016 0.468 ;
        RECT 1.572 0.54 1.764 0.612 ;
        RECT 1.692 0.396 1.764 0.612 ;
      LAYER V0 ;
        RECT 1.908 0.396 1.98 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 1.116 0.468 ;
        RECT 0.504 0.252 0.576 0.468 ;
        RECT 0.376 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 2.76 0.648 2.856 0.912 ;
        RECT 2.328 0.648 2.424 0.912 ;
        RECT 1.896 0.648 1.992 0.912 ;
        RECT 1.464 0.648 1.56 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.684 2.952 0.756 ;
        RECT 2.88 0.252 2.952 0.756 ;
        RECT 2.34 0.252 2.952 0.324 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.34 0.252 2.412 0.324 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.772 0.252 2.844 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.672 0.108 2.648 0.18 ;
      RECT 1.024 0.252 2 0.324 ;
      RECT 0.376 0.108 1.352 0.18 ;
  END
END NAND4xp75_ASAP7_6t_fix

MACRO NAND5xp2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND5xp2_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.576 0.18 ;
        RECT 0.288 0.108 0.36 0.504 ;
      LAYER V0 ;
        RECT 0.288 0.396 0.36 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.36 0.576 0.584 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 1.008 0.18 ;
        RECT 0.72 0.108 0.792 0.584 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.328 1.008 0.584 ;
      LAYER V0 ;
        RECT 0.936 0.38 1.008 0.452 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.52 1.44 0.728 ;
        RECT 1.152 0.108 1.44 0.18 ;
        RECT 1.152 0.52 1.44 0.592 ;
        RECT 1.152 0.108 1.224 0.592 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 1.136 0.756 ;
        RECT 0.072 0.212 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.232 0.144 0.304 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 1.044 0.684 1.116 0.756 ;
    END
  END Y
END NAND5xp2_ASAP7_6t_fix

MACRO NOR2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.148 0.54 0.296 0.612 ;
        RECT 0.148 0.108 0.296 0.18 ;
        RECT 0.148 0.108 0.22 0.612 ;
      LAYER V0 ;
        RECT 0.148 0.396 0.22 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1 0.54 1.224 0.612 ;
        RECT 1.152 0.108 1.224 0.612 ;
        RECT 0.676 0.396 1.224 0.468 ;
        RECT 1.076 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.54 0.9 0.612 ;
        RECT 0.396 0.108 0.9 0.18 ;
        RECT 0.396 0.108 0.468 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.252 0.468 0.324 ;
        RECT 0.828 0.54 0.9 0.612 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.684 1.116 0.756 ;
  END
END NOR2x1_ASAP7_6t_fix

MACRO NOR2x1p5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1p5_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 1.332 0.468 ;
        RECT 0.384 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.384 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 1.26 0.396 1.332 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 0.396 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.476 0.684 1.548 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.54 1.332 0.612 ;
      RECT 0.396 0.684 0.9 0.756 ;
  END
END NOR2x1p5_ASAP7_6t_fix

MACRO NOR2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.204 0.468 ;
        RECT 0.8 0.54 1.16 0.612 ;
        RECT 0.936 0.396 1.008 0.612 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.464 0.396 1.808 0.468 ;
        RECT 1.464 0.252 1.536 0.468 ;
        RECT 0.62 0.252 1.536 0.324 ;
        RECT 0.396 0.396 0.692 0.468 ;
        RECT 0.62 0.252 0.692 0.468 ;
      LAYER V0 ;
        RECT 0.396 0.396 0.468 0.468 ;
        RECT 1.692 0.396 1.764 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.54 2.088 0.612 ;
        RECT 2.016 0.108 2.088 0.612 ;
        RECT 0.072 0.108 2.088 0.18 ;
        RECT 0.072 0.54 0.468 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.54 0.468 0.612 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.54 1.764 0.612 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 2 0.756 ;
  END
END NOR2x2_ASAP7_6t_fix

MACRO NOR2xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp33_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.448 0.756 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.244 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.356 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.572 0.684 0.792 0.756 ;
        RECT 0.72 0.108 0.792 0.756 ;
        RECT 0.396 0.108 0.792 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.612 0.684 0.684 0.756 ;
    END
  END Y
END NOR2xp33_ASAP7_6t_fix

MACRO NOR2xp67_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2xp67_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.396 0.18 ;
        RECT 0.072 0.54 0.38 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.396 0.9 0.468 ;
        RECT 0.504 0.252 0.576 0.468 ;
        RECT 0.364 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.396 0.9 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.54 1.224 0.612 ;
        RECT 1.152 0.108 1.224 0.612 ;
        RECT 0.572 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 0.828 0.54 0.9 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 1.136 0.756 ;
  END
END NOR2xp67_ASAP7_6t_fix

MACRO NOR3x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.824 0.396 2.304 0.468 ;
        RECT 2.232 0.108 2.304 0.468 ;
        RECT 2.008 0.108 2.304 0.18 ;
      LAYER V0 ;
        RECT 1.908 0.396 1.98 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.128 0.252 1.352 0.324 ;
        RECT 0.936 0.396 1.2 0.468 ;
        RECT 1.128 0.252 1.2 0.468 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.684 0.18 ;
        RECT 0.072 0.54 0.22 0.612 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
        RECT 0.16 0.684 0.704 0.756 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
        RECT 0.6 0.54 0.696 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.54 2.216 0.612 ;
        RECT 0.808 0.108 1.764 0.18 ;
        RECT 1.512 0.108 1.584 0.612 ;
      LAYER V0 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.692 0.54 1.764 0.612 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.54 2.196 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.684 2 0.756 ;
      RECT 0.396 0.54 1.332 0.612 ;
  END
END NOR3x1_ASAP7_6t_fix

MACRO NOR3x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2_ASAP7_6t_fix 0 0 ;
  SIZE 4.32 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.904 0.396 3.148 0.468 ;
        RECT 2.904 0.252 2.976 0.468 ;
        RECT 1.132 0.252 2.976 0.324 ;
        RECT 0.928 0.396 1.204 0.468 ;
        RECT 1.132 0.252 1.204 0.468 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
        RECT 2.988 0.396 3.06 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.328 0.396 2.78 0.468 ;
      LAYER V0 ;
        RECT 2.124 0.396 2.196 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 4.32 0.9 ;
        RECT 1.672 0.684 2.648 0.756 ;
      LAYER LISD ;
        RECT 0 0.816 4.32 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 2.544 0.54 2.64 0.756 ;
        RECT 1.68 0.54 1.776 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 4.32 0.048 ;
        RECT 3.408 -0.048 3.504 0.324 ;
        RECT 2.976 -0.048 3.072 0.324 ;
        RECT 2.544 -0.048 2.64 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.616 0.54 4.248 0.612 ;
        RECT 4.176 0.108 4.248 0.612 ;
        RECT 0.528 0.108 4.248 0.18 ;
      LAYER V0 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.476 0.108 1.548 0.18 ;
        RECT 2.772 0.108 2.844 0.18 ;
        RECT 3.636 0.54 3.708 0.612 ;
        RECT 3.636 0.108 3.708 0.18 ;
        RECT 4.068 0.54 4.14 0.612 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.428 0.252 3.896 0.324 ;
      LAYER M1 ;
        RECT 3.724 0.252 3.888 0.324 ;
        RECT 3.552 0.396 3.796 0.468 ;
        RECT 3.724 0.252 3.796 0.468 ;
        RECT 0.528 0.396 0.684 0.468 ;
        RECT 0.528 0.252 0.6 0.468 ;
        RECT 0.436 0.252 0.6 0.324 ;
      LAYER V1 ;
        RECT 0.456 0.252 0.528 0.324 ;
        RECT 3.796 0.252 3.868 0.324 ;
      LAYER V0 ;
        RECT 0.612 0.396 0.684 0.468 ;
        RECT 3.636 0.396 3.708 0.468 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 2.968 0.684 3.944 0.756 ;
      RECT 1.044 0.54 3.296 0.612 ;
      RECT 0.376 0.684 1.352 0.756 ;
      RECT 0.18 0.54 0.684 0.612 ;
  END
END NOR3x2_ASAP7_6t_fix

MACRO NOR3xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.252 0.716 0.324 ;
        RECT 0.316 0.54 0.556 0.612 ;
        RECT 0.316 0.252 0.388 0.612 ;
      LAYER V0 ;
        RECT 0.316 0.396 0.388 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.344 0.684 0.952 0.756 ;
        RECT 0.88 0.396 0.952 0.756 ;
        RECT 0.512 0.396 0.952 0.468 ;
      LAYER V0 ;
        RECT 0.532 0.396 0.604 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 0.828 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.704 0.18 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.54 0.144 0.612 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
END NOR3xp33_ASAP7_6t_fix

MACRO NOR4xp25_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp25_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.224 0.612 ;
        RECT 0.936 0.252 1.224 0.324 ;
        RECT 0.936 0.252 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.684 0.968 0.756 ;
        RECT 0.72 0.252 0.792 0.756 ;
        RECT 0.572 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.336 0.396 0.596 0.468 ;
        RECT 0.336 0.684 0.576 0.756 ;
        RECT 0.336 0.396 0.408 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.36 0.324 ;
        RECT 0.072 0.684 0.236 0.756 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.208 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 0.16 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
END NOR4xp25_ASAP7_6t_fix

MACRO NOR4xp75_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4xp75_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.664 0.396 2.952 0.468 ;
        RECT 2.88 0.108 2.952 0.468 ;
        RECT 2.8 0.108 2.952 0.18 ;
      LAYER V0 ;
        RECT 2.772 0.396 2.844 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.728 0.396 2 0.468 ;
        RECT 1.728 0.252 1.8 0.468 ;
        RECT 1.512 0.252 1.8 0.324 ;
      LAYER V0 ;
        RECT 1.908 0.396 1.98 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.3 0.468 ;
        RECT 0.936 0.252 1.008 0.468 ;
        RECT 0.5 0.252 1.008 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 2.76 -0.048 2.856 0.216 ;
        RECT 2.328 -0.048 2.424 0.216 ;
        RECT 1.896 -0.048 1.992 0.216 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 1.032 -0.048 1.128 0.216 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 0.54 2.844 0.612 ;
        RECT 0.376 0.108 2.628 0.18 ;
        RECT 2.448 0.108 2.52 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.108 0.9 0.18 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.108 2.196 0.18 ;
        RECT 2.34 0.54 2.412 0.612 ;
        RECT 2.556 0.108 2.628 0.18 ;
        RECT 2.772 0.54 2.844 0.612 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.672 0.684 2.648 0.756 ;
      RECT 1.024 0.54 2 0.612 ;
      RECT 0.376 0.684 1.352 0.756 ;
  END
END NOR4xp75_ASAP7_6t_fix

MACRO NOR5xp2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR5xp2_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.252 0.452 0.324 ;
        RECT 0.288 0.252 0.36 0.584 ;
      LAYER V0 ;
        RECT 0.288 0.396 0.36 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.684 0.576 0.756 ;
        RECT 0.504 0.392 0.576 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.412 0.576 0.484 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.728 ;
        RECT 0.628 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.684 1.084 0.756 ;
        RECT 0.936 0.252 1.084 0.324 ;
        RECT 0.936 0.252 1.008 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.292 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 1.292 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.216 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 1.136 0.18 ;
        RECT 0.072 0.684 0.272 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.612 0.108 0.684 0.18 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
END NOR5xp2_ASAP7_6t_fix

MACRO O2A1O1Ixp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1Ixp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.656 0.54 0.876 0.612 ;
        RECT 0.804 0.396 0.876 0.612 ;
        RECT 0.3 0.396 0.876 0.468 ;
      LAYER V0 ;
        RECT 0.52 0.396 0.592 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.272 0.756 ;
        RECT 0.072 0.252 0.232 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.684 1.172 0.756 ;
        RECT 1.024 0.252 1.172 0.324 ;
        RECT 1.024 0.252 1.096 0.756 ;
      LAYER V0 ;
        RECT 1.024 0.396 1.096 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.684 1.656 0.756 ;
        RECT 1.584 0.252 1.656 0.756 ;
        RECT 1.348 0.396 1.656 0.468 ;
        RECT 1.424 0.252 1.656 0.324 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 0.816 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.108 1.568 0.18 ;
        RECT 0.356 0.252 0.88 0.324 ;
        RECT 0.808 0.108 0.88 0.324 ;
      LAYER V0 ;
        RECT 0.376 0.252 0.448 0.324 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.9 0.756 ;
      RECT 0.16 0.108 0.684 0.18 ;
  END
END O2A1O1Ixp33_ASAP7_6t_fix

MACRO O2A1O1Ixp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1Ixp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.464 ;
        RECT 0.288 0.252 1.008 0.324 ;
        RECT 0.288 0.108 0.36 0.324 ;
        RECT 0.072 0.108 0.36 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 0.936 0.392 1.008 0.464 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.396 0.724 0.468 ;
        RECT 0.072 0.684 0.288 0.756 ;
        RECT 0.216 0.396 0.288 0.756 ;
      LAYER V0 ;
        RECT 0.612 0.396 0.684 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.036 0.54 1.224 0.612 ;
        RECT 1.152 0.28 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.392 1.224 0.464 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.324 0.54 1.472 0.612 ;
        RECT 1.368 0.28 1.44 0.612 ;
      LAYER V0 ;
        RECT 1.368 0.392 1.44 0.464 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.108 1.656 0.704 ;
        RECT 1.26 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.584 0.612 1.656 0.684 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.504 0.684 1.332 0.756 ;
      RECT 0.612 0.108 1.116 0.18 ;
      RECT 0.396 0.54 0.872 0.612 ;
  END
END O2A1O1Ixp5_ASAP7_6t_fix

MACRO OA211x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.412 0.54 0.58 0.612 ;
        RECT 0.508 0.396 0.58 0.612 ;
      LAYER V0 ;
        RECT 0.508 0.468 0.58 0.54 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.108 1.016 0.18 ;
        RECT 0.72 0.468 0.864 0.54 ;
        RECT 0.792 0.108 0.864 0.54 ;
      LAYER V0 ;
        RECT 0.72 0.468 0.792 0.54 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.14 0.324 ;
        RECT 0.936 0.54 1.084 0.612 ;
        RECT 0.936 0.252 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.108 1.44 0.728 ;
        RECT 1.14 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 1.368 0.204 1.44 0.276 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.216 0.684 1.292 0.756 ;
      RECT 1.22 0.396 1.292 0.756 ;
      RECT 0.216 0.252 0.288 0.756 ;
      RECT 0.216 0.252 0.44 0.324 ;
      RECT 0.18 0.108 0.684 0.18 ;
  END
END OA211x1_ASAP7_6t_fix

MACRO OA211x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.54 0.576 0.612 ;
        RECT 0.504 0.424 0.576 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.468 0.576 0.54 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.38 0.468 ;
        RECT 0.072 0.252 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.22 0.396 0.292 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.56 ;
        RECT 0.632 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.468 0.792 0.54 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.008 0.552 ;
        RECT 0.828 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.24 0.108 1.656 0.18 ;
        RECT 1.296 0.612 1.368 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.296 0.612 1.368 0.684 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.684 1.164 0.756 ;
      RECT 1.092 0.252 1.164 0.756 ;
      RECT 1.092 0.396 1.312 0.468 ;
      RECT 1.092 0.252 1.344 0.324 ;
      RECT 0.18 0.108 0.704 0.18 ;
      RECT 0.34 0.252 0.508 0.324 ;
    LAYER M2 ;
      RECT 0.376 0.252 1.24 0.324 ;
    LAYER V1 ;
      RECT 1.168 0.252 1.24 0.324 ;
      RECT 0.396 0.252 0.468 0.324 ;
  END
END OA211x2_ASAP7_6t_fix

MACRO OA21x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.384 0.396 0.624 0.468 ;
        RECT 0.384 0.54 0.604 0.612 ;
        RECT 0.384 0.396 0.456 0.612 ;
      LAYER V0 ;
        RECT 0.532 0.396 0.604 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.748 0.396 1.12 0.468 ;
        RECT 1.048 0.252 1.12 0.468 ;
        RECT 0.9 0.252 1.12 0.324 ;
      LAYER V0 ;
        RECT 0.748 0.396 0.82 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 1.008 0.108 1.44 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.232 0.684 0.9 0.756 ;
      RECT 0.828 0.54 0.9 0.756 ;
      RECT 0.232 0.252 0.304 0.756 ;
      RECT 0.828 0.54 1.28 0.612 ;
      RECT 1.208 0.38 1.28 0.612 ;
      RECT 0.232 0.252 0.516 0.324 ;
      RECT 0.18 0.108 0.684 0.18 ;
  END
END OA21x2_ASAP7_6t_fix

MACRO OA221x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221x1_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.568 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.572 0.396 0.792 0.468 ;
        RECT 0.244 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.612 0.396 0.684 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.236 0.612 ;
        RECT 0.936 0.396 1.224 0.468 ;
        RECT 0.936 0.396 1.008 0.612 ;
      LAYER V0 ;
        RECT 1.044 0.396 1.116 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.188 0.54 2.52 0.612 ;
        RECT 2.448 0.396 2.52 0.612 ;
        RECT 2.188 0.396 2.52 0.468 ;
      LAYER V0 ;
        RECT 2.34 0.396 2.412 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.364 0.54 2.088 0.612 ;
        RECT 2.016 0.396 2.088 0.612 ;
        RECT 1.364 0.396 2.088 0.468 ;
      LAYER V0 ;
        RECT 1.908 0.396 1.98 0.468 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.664 0.54 2.996 0.612 ;
        RECT 2.664 0.396 2.996 0.468 ;
        RECT 2.664 0.396 2.736 0.612 ;
      LAYER V0 ;
        RECT 2.772 0.396 2.844 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.544 0.54 2.64 0.912 ;
        RECT 2.328 0.54 2.64 0.756 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.616 0.828 0.688 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.36 0.18 ;
        RECT 0.072 0.684 0.252 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 0.18 0.108 0.252 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 3.168 0.756 ;
      RECT 3.096 0.252 3.168 0.756 ;
      RECT 0.396 0.396 0.468 0.756 ;
      RECT 0.244 0.396 0.468 0.468 ;
      RECT 2.556 0.252 3.168 0.324 ;
      RECT 1.26 0.252 2.412 0.324 ;
      RECT 1.26 0.108 1.332 0.324 ;
      RECT 0.576 0.108 1.332 0.18 ;
      RECT 1.692 0.108 3.08 0.18 ;
  END
END OA221x1_ASAP7_6t_fix

MACRO OA221x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221x2_ASAP7_6t_fix 0 0 ;
  SIZE 3.456 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.864 0.396 1.028 0.468 ;
        RECT 0.864 0.252 0.936 0.468 ;
        RECT 0.284 0.252 0.936 0.324 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.54 1.668 0.612 ;
        RECT 1.368 0.252 1.44 0.612 ;
        RECT 1.156 0.252 1.44 0.324 ;
      LAYER V0 ;
        RECT 1.368 0.404 1.44 0.476 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 0.54 2.704 0.612 ;
        RECT 2.52 0.404 2.592 0.612 ;
        RECT 2.408 0.404 2.592 0.476 ;
      LAYER V0 ;
        RECT 2.448 0.404 2.52 0.476 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.944 0.4 2.128 0.472 ;
        RECT 1.792 0.54 2.016 0.612 ;
        RECT 1.944 0.4 2.016 0.612 ;
      LAYER V0 ;
        RECT 2.016 0.4 2.088 0.472 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.948 0.54 3.168 0.612 ;
        RECT 3.096 0.396 3.168 0.612 ;
        RECT 2.792 0.396 3.168 0.468 ;
      LAYER V0 ;
        RECT 2.988 0.396 3.06 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.456 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.456 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.544 0.54 2.856 0.756 ;
        RECT 2.544 0.54 2.64 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.832 0.828 0.904 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.456 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.684 0.468 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.576 0.684 3.384 0.756 ;
      RECT 3.312 0.252 3.384 0.756 ;
      RECT 0.576 0.396 0.648 0.756 ;
      RECT 0.484 0.396 0.648 0.468 ;
      RECT 2.988 0.252 3.384 0.324 ;
      RECT 1.656 0.252 2.652 0.324 ;
      RECT 1.656 0.108 1.728 0.324 ;
      RECT 0.828 0.108 1.728 0.18 ;
      RECT 1.908 0.108 3.296 0.18 ;
  END
END OA221x2_ASAP7_6t_fix

MACRO OA222x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.396 0.5 0.468 ;
        RECT 0.216 0.54 0.492 0.612 ;
        RECT 0.216 0.396 0.288 0.612 ;
      LAYER V0 ;
        RECT 0.292 0.396 0.364 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.54 0.792 0.612 ;
        RECT 0.72 0.324 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.348 0.54 1.656 0.612 ;
        RECT 1.584 0.396 1.656 0.612 ;
        RECT 1.348 0.396 1.656 0.468 ;
      LAYER V0 ;
        RECT 1.44 0.396 1.512 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.408 1.196 0.48 ;
        RECT 0.932 0.54 1.08 0.612 ;
        RECT 1.008 0.252 1.08 0.612 ;
        RECT 0.932 0.252 1.08 0.324 ;
      LAYER V0 ;
        RECT 1.124 0.408 1.196 0.48 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.54 2.172 0.612 ;
        RECT 1.8 0.396 1.872 0.612 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 0.108 2.54 0.18 ;
        RECT 1.992 0.252 2.392 0.324 ;
        RECT 2.32 0.108 2.392 0.324 ;
        RECT 2.232 0.252 2.304 0.46 ;
      LAYER V0 ;
        RECT 2.232 0.388 2.304 0.46 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.556 0.684 2.736 0.756 ;
        RECT 2.664 0.252 2.736 0.756 ;
      LAYER V0 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.664 0.252 2.736 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.684 2.424 0.756 ;
      RECT 2.352 0.548 2.424 0.756 ;
      RECT 0.072 0.252 0.144 0.756 ;
      RECT 2.352 0.548 2.504 0.62 ;
      RECT 2.432 0.4 2.504 0.62 ;
      RECT 0.072 0.252 0.544 0.324 ;
      RECT 1.26 0.252 1.764 0.324 ;
      RECT 1.692 0.108 1.764 0.324 ;
      RECT 1.692 0.108 2.196 0.18 ;
      RECT 0.18 0.108 1.568 0.18 ;
  END
END OA222x1_ASAP7_6t_fix

MACRO OA222x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222x2_ASAP7_6t_fix 0 0 ;
  SIZE 3.024 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.612 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.54 1.744 0.612 ;
        RECT 1.584 0.396 1.656 0.612 ;
        RECT 1.132 0.396 1.656 0.468 ;
      LAYER V0 ;
        RECT 1.44 0.396 1.512 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.44 0.612 ;
        RECT 0.936 0.252 1.156 0.324 ;
        RECT 0.936 0.252 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.844 0.252 2.124 0.324 ;
        RECT 1.672 0.684 1.916 0.756 ;
        RECT 1.844 0.252 1.916 0.756 ;
      LAYER V0 ;
        RECT 1.844 0.396 1.916 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.252 2.736 0.324 ;
        RECT 2.016 0.54 2.304 0.612 ;
        RECT 2.232 0.252 2.304 0.612 ;
      LAYER V0 ;
        RECT 2.232 0.408 2.304 0.48 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.024 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.024 0.912 ;
        RECT 2.76 0.54 2.856 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 0.6 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.024 0.048 ;
        RECT 2.76 -0.048 2.856 0.324 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.556 0.684 2.952 0.756 ;
        RECT 2.88 0.108 2.952 0.756 ;
        RECT 2.536 0.108 2.952 0.18 ;
      LAYER V0 ;
        RECT 2.556 0.684 2.628 0.756 ;
        RECT 2.556 0.108 2.628 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.124 0.684 2.456 0.756 ;
      RECT 2.384 0.396 2.456 0.756 ;
      RECT 2.384 0.396 2.648 0.468 ;
      RECT 1.28 0.252 1.744 0.324 ;
      RECT 1.672 0.108 1.744 0.324 ;
      RECT 1.672 0.108 2.304 0.18 ;
      RECT 0.324 0.684 1.548 0.756 ;
      RECT 0.324 0.252 0.396 0.756 ;
      RECT 0.324 0.252 0.488 0.324 ;
      RECT 0.18 0.108 1.548 0.18 ;
  END
END OA222x2_ASAP7_6t_fix

MACRO OA22x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.576 0.396 1.192 0.468 ;
        RECT 0.072 0.684 0.648 0.756 ;
        RECT 0.576 0.396 0.648 0.756 ;
        RECT 0.072 0.244 0.144 0.756 ;
      LAYER V0 ;
        RECT 1.08 0.396 1.152 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.932 0.54 1.44 0.612 ;
        RECT 1.368 0.408 1.44 0.612 ;
      LAYER V0 ;
        RECT 1.368 0.408 1.44 0.48 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.936 0.684 2.088 0.756 ;
        RECT 2.016 0.252 2.088 0.756 ;
        RECT 1.936 0.252 2.088 0.324 ;
      LAYER V0 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.54 1.736 0.612 ;
        RECT 1.584 0.252 1.732 0.324 ;
        RECT 1.584 0.252 1.656 0.612 ;
      LAYER V0 ;
        RECT 1.584 0.4 1.656 0.472 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.54 0.468 0.612 ;
        RECT 0.288 0.108 0.468 0.18 ;
        RECT 0.288 0.108 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.396 0.54 0.468 0.612 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.108 2 0.18 ;
      RECT 0.828 0.684 1.624 0.756 ;
      RECT 0.828 0.252 1.308 0.324 ;
  END
END OA22x2_ASAP7_6t_fix

MACRO OA31x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31x2_ASAP7_6t_fix 0 0 ;
  SIZE 3.24 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.312 0.612 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.396 0.832 0.468 ;
        RECT 0.432 0.54 0.692 0.612 ;
        RECT 0.432 0.396 0.504 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.328 0.396 1.804 0.468 ;
        RECT 1.328 0.252 1.4 0.468 ;
        RECT 1.252 0.252 1.4 0.324 ;
      LAYER V0 ;
        RECT 1.692 0.396 1.764 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.592 0.54 2.976 0.612 ;
        RECT 2.592 0.252 2.976 0.324 ;
        RECT 2.592 0.252 2.664 0.612 ;
        RECT 1.996 0.396 2.664 0.468 ;
      LAYER V0 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 3.24 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 3.24 0.912 ;
        RECT 2.976 0.54 3.072 0.912 ;
        RECT 2.544 0.54 2.64 0.912 ;
        RECT 2.112 0.648 2.208 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 3.24 0.048 ;
        RECT 2.976 -0.048 3.072 0.324 ;
        RECT 2.544 -0.048 2.64 0.324 ;
        RECT 2.112 -0.048 2.208 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.752 0.684 3.168 0.756 ;
        RECT 3.096 0.108 3.168 0.756 ;
        RECT 2.752 0.108 3.168 0.18 ;
      LAYER V0 ;
        RECT 2.772 0.684 2.844 0.756 ;
        RECT 2.772 0.108 2.844 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.268 0.684 1.784 0.756 ;
      RECT 1.268 0.54 1.34 0.756 ;
      RECT 0.832 0.54 1.34 0.612 ;
      RECT 0.632 0.252 1.116 0.324 ;
      RECT 0.632 0.108 0.704 0.324 ;
      RECT 0.072 0.108 0.704 0.18 ;
      RECT 1.524 0.252 2.444 0.324 ;
      RECT 1.476 0.54 2.444 0.612 ;
      RECT 0.828 0.108 2 0.18 ;
      RECT 0.16 0.684 1.136 0.756 ;
  END
END OA31x2_ASAP7_6t_fix

MACRO OA331x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.836 0.684 0.984 0.756 ;
        RECT 0.912 0.384 0.984 0.756 ;
      LAYER V0 ;
        RECT 0.912 0.408 0.984 0.48 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.676 0.252 0.824 0.324 ;
        RECT 0.644 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.4 0.792 0.472 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.464 ;
        RECT 0.416 0.252 0.576 0.324 ;
        RECT 0.416 0.108 0.488 0.324 ;
        RECT 0.28 0.108 0.488 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.392 0.576 0.464 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.064 0.684 1.212 0.756 ;
        RECT 1.064 0.396 1.212 0.468 ;
        RECT 1.064 0.396 1.136 0.756 ;
      LAYER V0 ;
        RECT 1.14 0.396 1.212 0.468 ;
    END
  END B1
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.612 0.252 1.88 0.324 ;
        RECT 1.436 0.54 1.684 0.612 ;
        RECT 1.612 0.252 1.684 0.612 ;
      LAYER V0 ;
        RECT 1.612 0.408 1.684 0.48 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.856 0.396 2.088 0.468 ;
        RECT 2.016 0.108 2.088 0.468 ;
        RECT 1.936 0.108 2.088 0.18 ;
      LAYER V0 ;
        RECT 1.856 0.396 1.928 0.468 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.244 0.144 0.62 ;
      LAYER V0 ;
        RECT 0.072 0.412 0.144 0.484 ;
    END
  END Y
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.368 0.396 1.572 0.468 ;
      LAYER M1 ;
        RECT 1.34 0.396 1.488 0.468 ;
      LAYER V1 ;
        RECT 1.368 0.396 1.44 0.468 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B2
  OBS
    LAYER M1 ;
      RECT 1.044 0.252 1.512 0.324 ;
      RECT 1.044 0.108 1.116 0.324 ;
      RECT 0.612 0.108 1.116 0.18 ;
      RECT 0.372 0.684 0.684 0.756 ;
      RECT 0.372 0.532 0.444 0.756 ;
      RECT 0.288 0.532 0.444 0.604 ;
      RECT 0.288 0.412 0.36 0.604 ;
      RECT 1.476 0.684 2 0.756 ;
      RECT 1.26 0.108 1.788 0.18 ;
  END
END OA331x1_ASAP7_6t_fix

MACRO OA331x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 -1.104 ;
  FOREIGN OA331x2_ASAP7_6t_fix 0 1.104 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.072 1.5 1.24 1.572 ;
      LAYER M1 ;
        RECT 1.128 1.488 1.2 1.66 ;
        RECT 0.064 1.712 0.212 1.86 ;
        RECT 0.064 1.212 0.212 1.428 ;
        RECT 0.092 1.212 0.164 1.86 ;
      LAYER V1 ;
        RECT 0.092 1.5 0.164 1.572 ;
        RECT 1.128 1.5 1.2 1.572 ;
      LAYER V0 ;
        RECT 1.128 1.512 1.2 1.584 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.892 1.356 1.04 1.428 ;
        RECT 0.876 1.644 1.024 1.716 ;
        RECT 0.936 1.356 1.008 1.716 ;
      LAYER V0 ;
        RECT 0.936 1.504 1.008 1.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 1.356 0.792 1.568 ;
        RECT 0.632 1.356 0.792 1.428 ;
        RECT 0.632 1.212 0.704 1.428 ;
        RECT 0.352 1.212 0.704 1.284 ;
      LAYER V0 ;
        RECT 0.72 1.496 0.792 1.568 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.28 1.712 1.428 1.86 ;
        RECT 1.28 1.512 1.428 1.584 ;
        RECT 1.28 1.512 1.352 1.86 ;
      LAYER V0 ;
        RECT 1.356 1.512 1.428 1.584 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.632 1.788 1.78 1.86 ;
        RECT 1.632 1.512 1.704 1.86 ;
        RECT 1.556 1.512 1.704 1.584 ;
      LAYER V0 ;
        RECT 1.556 1.512 1.628 1.584 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.828 1.644 2.244 1.716 ;
        RECT 1.828 1.492 1.9 1.716 ;
      LAYER V0 ;
        RECT 1.828 1.512 1.9 1.584 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.072 1.5 2.304 1.572 ;
        RECT 2.156 1.212 2.304 1.572 ;
      LAYER V0 ;
        RECT 2.072 1.5 2.144 1.572 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.932 2.376 2.004 ;
      LAYER LISD ;
        RECT 0 1.92 2.376 2.016 ;
        RECT 1.896 1.644 1.992 2.016 ;
        RECT 0.6 1.644 0.696 2.016 ;
        RECT 0.168 1.644 0.264 2.016 ;
      LAYER V0 ;
        RECT 0.18 1.932 0.252 2.004 ;
        RECT 0.396 1.932 0.468 2.004 ;
        RECT 0.612 1.932 0.684 2.004 ;
        RECT 0.828 1.932 0.9 2.004 ;
        RECT 1.044 1.932 1.116 2.004 ;
        RECT 1.26 1.932 1.332 2.004 ;
        RECT 1.476 1.932 1.548 2.004 ;
        RECT 1.692 1.932 1.764 2.004 ;
        RECT 1.908 1.932 1.98 2.004 ;
        RECT 2.124 1.932 2.196 2.004 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.068 2.376 1.14 ;
      LAYER LISD ;
        RECT 0 1.056 2.376 1.152 ;
        RECT 1.032 1.056 1.128 1.428 ;
        RECT 0.6 1.056 0.696 1.428 ;
        RECT 0.168 1.056 0.264 1.428 ;
      LAYER V0 ;
        RECT 0.18 1.068 0.252 1.14 ;
        RECT 0.396 1.068 0.468 1.14 ;
        RECT 0.612 1.068 0.684 1.14 ;
        RECT 0.828 1.068 0.9 1.14 ;
        RECT 1.044 1.068 1.116 1.14 ;
        RECT 1.26 1.068 1.332 1.14 ;
        RECT 1.476 1.068 1.548 1.14 ;
        RECT 1.692 1.068 1.764 1.14 ;
        RECT 1.908 1.068 1.98 1.14 ;
        RECT 2.124 1.068 2.196 1.14 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 1.788 0.468 1.86 ;
        RECT 0.288 1.356 0.456 1.428 ;
        RECT 0.288 1.356 0.36 1.86 ;
      LAYER V0 ;
        RECT 0.36 1.356 0.432 1.428 ;
        RECT 0.396 1.788 0.468 1.86 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.26 1.356 1.78 1.428 ;
      RECT 1.26 1.212 1.332 1.428 ;
      RECT 0.828 1.212 1.332 1.284 ;
      RECT 0.588 1.788 0.74 1.86 ;
      RECT 0.588 1.636 0.66 1.86 ;
      RECT 0.504 1.636 0.66 1.708 ;
      RECT 0.504 1.516 0.576 1.708 ;
      RECT 2.068 1.788 2.216 1.86 ;
      RECT 1.476 1.212 2.004 1.284 ;
      RECT 1.012 1.788 1.16 1.86 ;
    LAYER M2 ;
      RECT 0.64 1.788 2.216 1.86 ;
    LAYER V1 ;
      RECT 2.124 1.788 2.196 1.86 ;
      RECT 1.044 1.788 1.116 1.86 ;
      RECT 0.66 1.788 0.732 1.86 ;
  END
END OA331x2_ASAP7_6t_fix

MACRO OA332x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.408 0.98 0.728 ;
      LAYER V0 ;
        RECT 0.908 0.408 0.98 0.48 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.868 0.324 ;
        RECT 0.4 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.4 0.792 0.472 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.396 0.648 0.468 ;
        RECT 0.576 0.252 0.648 0.468 ;
        RECT 0.316 0.252 0.648 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.052 0.396 1.2 0.468 ;
        RECT 1.052 0.396 1.124 0.728 ;
      LAYER V0 ;
        RECT 1.128 0.396 1.2 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.416 0.408 1.488 0.728 ;
        RECT 1.34 0.408 1.488 0.48 ;
      LAYER V0 ;
        RECT 1.34 0.408 1.412 0.48 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.608 0.388 1.68 0.688 ;
      LAYER V0 ;
        RECT 1.608 0.408 1.68 0.48 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.932 0.396 2.14 0.468 ;
        RECT 1.932 0.396 2.004 0.724 ;
      LAYER V0 ;
        RECT 2.068 0.396 2.14 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.788 0.388 1.86 0.688 ;
      LAYER V0 ;
        RECT 1.788 0.408 1.86 0.48 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.108 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.408 0.144 0.48 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.164 0.684 2.312 0.756 ;
      RECT 2.24 0.252 2.312 0.756 ;
      RECT 1.908 0.252 2.312 0.324 ;
      RECT 1.044 0.252 1.56 0.324 ;
      RECT 1.044 0.108 1.116 0.324 ;
      RECT 0.612 0.108 1.116 0.18 ;
      RECT 0.228 0.684 0.808 0.756 ;
      RECT 0.228 0.408 0.3 0.756 ;
      RECT 1.26 0.108 2.224 0.18 ;
    LAYER M2 ;
      RECT 0.708 0.684 2.296 0.756 ;
    LAYER V1 ;
      RECT 2.204 0.684 2.276 0.756 ;
      RECT 0.728 0.684 0.8 0.756 ;
  END
END OA332x1_ASAP7_6t_fix

MACRO OA332x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.54 1.224 0.612 ;
        RECT 1.152 0.408 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.408 1.224 0.48 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.252 1.096 0.324 ;
        RECT 0.908 0.252 0.98 0.488 ;
      LAYER V0 ;
        RECT 0.908 0.396 0.98 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.62 0.54 0.768 0.612 ;
        RECT 0.696 0.252 0.768 0.612 ;
        RECT 0.36 0.252 0.768 0.324 ;
        RECT 0.36 0.396 0.58 0.468 ;
        RECT 0.36 0.252 0.432 0.468 ;
      LAYER V0 ;
        RECT 0.696 0.396 0.768 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.684 1.444 0.756 ;
        RECT 1.296 0.396 1.444 0.468 ;
        RECT 1.296 0.396 1.368 0.756 ;
      LAYER V0 ;
        RECT 1.372 0.396 1.444 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.588 0.684 1.752 0.756 ;
        RECT 1.68 0.428 1.752 0.756 ;
        RECT 1.568 0.428 1.752 0.5 ;
      LAYER V0 ;
        RECT 1.588 0.428 1.66 0.5 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.824 0.388 1.896 0.688 ;
      LAYER V0 ;
        RECT 1.824 0.408 1.896 0.48 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.208 0.408 2.356 0.48 ;
        RECT 2.208 0.408 2.28 0.728 ;
      LAYER V0 ;
        RECT 2.284 0.408 2.356 0.48 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.004 0.388 2.076 0.688 ;
      LAYER V0 ;
        RECT 2.004 0.408 2.076 0.48 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.108 0.468 0.18 ;
        RECT 0.216 0.54 0.44 0.612 ;
        RECT 0.216 0.108 0.288 0.612 ;
      LAYER V0 ;
        RECT 0.348 0.54 0.42 0.612 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.38 0.684 2.528 0.756 ;
      RECT 2.456 0.252 2.528 0.756 ;
      RECT 2.124 0.252 2.528 0.324 ;
      RECT 1.26 0.252 1.776 0.324 ;
      RECT 1.26 0.108 1.332 0.324 ;
      RECT 0.704 0.108 1.332 0.18 ;
      RECT 0.072 0.684 0.92 0.756 ;
      RECT 0.072 0.396 0.144 0.756 ;
      RECT 1.476 0.108 2.44 0.18 ;
    LAYER M2 ;
      RECT 0.808 0.684 2.512 0.756 ;
    LAYER V1 ;
      RECT 2.42 0.684 2.492 0.756 ;
      RECT 0.828 0.684 0.9 0.756 ;
  END
END OA332x2_ASAP7_6t_fix

MACRO OA333x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.18 0.684 2.528 0.756 ;
        RECT 2.456 0.396 2.528 0.756 ;
        RECT 2.296 0.396 2.528 0.468 ;
      LAYER V0 ;
        RECT 2.296 0.396 2.368 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.952 0.54 2.296 0.612 ;
        RECT 1.952 0.396 2.172 0.468 ;
        RECT 1.952 0.396 2.024 0.612 ;
      LAYER V0 ;
        RECT 2.024 0.396 2.104 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.792 0.396 1.864 0.612 ;
      LAYER V0 ;
        RECT 1.792 0.396 1.864 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.052 0.396 1.2 0.468 ;
        RECT 1.052 0.396 1.124 0.544 ;
      LAYER V0 ;
        RECT 1.128 0.396 1.2 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.352 0.608 1.512 0.756 ;
        RECT 1.416 0.396 1.488 0.756 ;
        RECT 1.34 0.396 1.488 0.468 ;
      LAYER V0 ;
        RECT 1.34 0.396 1.412 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.612 0.388 1.684 0.728 ;
      LAYER V0 ;
        RECT 1.612 0.408 1.684 0.48 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.492 0.684 0.98 0.756 ;
        RECT 0.908 0.408 0.98 0.756 ;
        RECT 0.492 0.54 0.564 0.756 ;
        RECT 0.4 0.54 0.564 0.612 ;
      LAYER V0 ;
        RECT 0.908 0.408 0.98 0.48 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.54 0.836 0.612 ;
        RECT 0.72 0.464 0.836 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.532 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.392 0.792 0.464 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.396 0.58 0.468 ;
        RECT 0.36 0.108 0.432 0.468 ;
        RECT 0.244 0.108 0.432 0.18 ;
      LAYER V0 ;
        RECT 0.476 0.396 0.548 0.468 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.136 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.252 0.144 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.908 0.252 2.52 0.324 ;
      RECT 1.908 0.16 1.98 0.324 ;
      RECT 1.044 0.252 1.54 0.324 ;
      RECT 1.044 0.108 1.116 0.324 ;
      RECT 0.612 0.108 1.116 0.18 ;
      RECT 0.216 0.684 0.364 0.756 ;
      RECT 0.216 0.408 0.288 0.756 ;
      RECT 2.124 0.108 2.276 0.18 ;
      RECT 1.908 0.684 2.056 0.756 ;
      RECT 1.26 0.108 1.764 0.18 ;
      RECT 1.08 0.684 1.24 0.756 ;
    LAYER M2 ;
      RECT 1.684 0.108 2.224 0.18 ;
      RECT 0.264 0.684 2.008 0.756 ;
    LAYER V1 ;
      RECT 2.132 0.108 2.204 0.18 ;
      RECT 1.916 0.684 1.988 0.756 ;
      RECT 1.684 0.108 1.756 0.18 ;
      RECT 1.124 0.684 1.196 0.756 ;
      RECT 0.284 0.684 0.356 0.756 ;
  END
END OA333x1_ASAP7_6t_fix

MACRO OA333x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.596 0.608 2.744 0.756 ;
        RECT 2.672 0.396 2.744 0.756 ;
        RECT 2.444 0.396 2.744 0.468 ;
      LAYER V0 ;
        RECT 2.444 0.396 2.516 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.168 0.408 2.32 0.48 ;
        RECT 2.168 0.408 2.24 0.728 ;
      LAYER V0 ;
        RECT 2.24 0.408 2.32 0.48 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.008 0.408 2.08 0.728 ;
      LAYER V0 ;
        RECT 2.008 0.408 2.08 0.48 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.268 0.396 1.416 0.468 ;
        RECT 1.268 0.396 1.34 0.544 ;
      LAYER V0 ;
        RECT 1.344 0.396 1.416 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.568 0.608 1.728 0.756 ;
        RECT 1.632 0.396 1.704 0.756 ;
        RECT 1.556 0.396 1.704 0.468 ;
      LAYER V0 ;
        RECT 1.556 0.396 1.628 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.828 0.388 1.9 0.728 ;
      LAYER V0 ;
        RECT 1.828 0.408 1.9 0.48 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.048 0.684 1.196 0.756 ;
        RECT 1.124 0.408 1.196 0.756 ;
      LAYER V0 ;
        RECT 1.124 0.408 1.196 0.48 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.892 0.252 1.04 0.324 ;
        RECT 0.86 0.536 1.008 0.608 ;
        RECT 0.936 0.252 1.008 0.608 ;
        RECT 0.784 0.684 0.932 0.756 ;
        RECT 0.86 0.536 0.932 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.452 ;
        RECT 0.632 0.252 0.792 0.324 ;
        RECT 0.632 0.108 0.704 0.324 ;
        RECT 0.284 0.108 0.704 0.18 ;
      LAYER V0 ;
        RECT 0.72 0.38 0.792 0.452 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.32 0.684 0.468 0.756 ;
        RECT 0.068 0.252 0.468 0.324 ;
        RECT 0.32 0.252 0.392 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.252 0.468 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.124 0.252 2.736 0.324 ;
      RECT 2.124 0.18 2.196 0.324 ;
      RECT 1.26 0.252 1.756 0.324 ;
      RECT 1.26 0.108 1.332 0.324 ;
      RECT 0.828 0.108 1.332 0.18 ;
      RECT 0.068 0.684 0.216 0.756 ;
      RECT 0.068 0.396 0.14 0.756 ;
      RECT 0.068 0.396 0.216 0.468 ;
      RECT 2.34 0.108 2.492 0.18 ;
      RECT 2.34 0.684 2.488 0.756 ;
      RECT 1.476 0.108 1.98 0.18 ;
      RECT 1.296 0.684 1.456 0.756 ;
    LAYER M2 ;
      RECT 1.9 0.108 2.484 0.18 ;
      RECT 0.072 0.684 2.44 0.756 ;
    LAYER V1 ;
      RECT 2.412 0.108 2.484 0.18 ;
      RECT 2.348 0.684 2.42 0.756 ;
      RECT 1.9 0.108 1.972 0.18 ;
      RECT 1.34 0.684 1.412 0.756 ;
      RECT 0.092 0.684 0.164 0.756 ;
  END
END OA333x2_ASAP7_6t_fix

MACRO OA33x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.54 ;
        RECT 0.384 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.892 0.252 1.04 0.324 ;
        RECT 0.936 0.252 1.008 0.552 ;
      LAYER V0 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 0.684 1.22 0.756 ;
        RECT 1.148 0.356 1.22 0.756 ;
      LAYER V0 ;
        RECT 1.148 0.396 1.22 0.468 ;
    END
  END A3
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 0.408 1.672 0.48 ;
        RECT 1.44 0.684 1.592 0.756 ;
        RECT 1.52 0.408 1.592 0.756 ;
      LAYER V0 ;
        RECT 1.592 0.408 1.672 0.48 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.34 0.28 1.412 0.56 ;
      LAYER V0 ;
        RECT 1.34 0.408 1.412 0.48 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.684 0.468 0.756 ;
        RECT 0.396 0.54 0.468 0.756 ;
        RECT 0.248 0.54 0.468 0.612 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.612 0.468 0.684 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.66 0.396 2.092 0.468 ;
      LAYER M1 ;
        RECT 1.872 0.396 1.944 0.572 ;
        RECT 1.796 0.396 1.944 0.468 ;
      LAYER V1 ;
        RECT 1.804 0.396 1.876 0.468 ;
      LAYER V0 ;
        RECT 1.796 0.396 1.868 0.468 ;
    END
  END B1
  OBS
    LAYER M1 ;
      RECT 1.692 0.684 2.088 0.756 ;
      RECT 2.016 0.252 2.088 0.756 ;
      RECT 1.484 0.252 2.088 0.324 ;
      RECT 1.484 0.16 1.556 0.324 ;
      RECT 0.576 0.684 0.9 0.756 ;
      RECT 0.576 0.396 0.648 0.756 ;
      RECT 0.388 0.396 0.648 0.468 ;
      RECT 1.692 0.108 1.844 0.18 ;
      RECT 0.792 0.108 1.332 0.18 ;
    LAYER M2 ;
      RECT 1.252 0.108 1.836 0.18 ;
    LAYER V1 ;
      RECT 1.764 0.108 1.836 0.18 ;
      RECT 1.252 0.108 1.324 0.18 ;
  END
END OA33x2_ASAP7_6t_fix

MACRO OAI211x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.484 0.396 0.812 0.468 ;
      LAYER V0 ;
        RECT 0.612 0.396 0.684 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.54 1.008 0.612 ;
        RECT 0.936 0.424 1.008 0.612 ;
        RECT 0.288 0.424 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.288 0.464 0.36 0.536 ;
        RECT 0.936 0.468 1.008 0.54 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.252 1.952 0.324 ;
        RECT 1.152 0.54 1.872 0.612 ;
        RECT 1.8 0.252 1.872 0.612 ;
        RECT 1.152 0.468 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.468 1.224 0.54 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.656 0.468 ;
        RECT 1.368 0.252 1.44 0.468 ;
        RECT 1.256 0.252 1.44 0.324 ;
      LAYER V0 ;
        RECT 1.468 0.396 1.54 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.68 0.648 1.776 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 1.98 0.756 ;
        RECT 0.072 0.252 0.9 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.448 0.144 0.52 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.252 0.468 0.324 ;
        RECT 0.828 0.252 0.9 0.324 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.908 0.684 1.98 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.98 0.18 ;
  END
END OAI211x1_ASAP7_6t_fix

MACRO OAI211xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.724 0.54 0.992 0.612 ;
        RECT 0.92 0.108 0.992 0.612 ;
        RECT 0.504 0.396 0.992 0.468 ;
        RECT 0.808 0.108 0.992 0.18 ;
      LAYER V0 ;
        RECT 0.576 0.396 0.648 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.224 0.756 ;
        RECT 0.072 0.252 0.224 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.54 1.388 0.612 ;
        RECT 1.08 0.108 1.244 0.18 ;
        RECT 1.08 0.108 1.152 0.612 ;
      LAYER V0 ;
        RECT 1.08 0.396 1.152 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.368 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.648 1.56 0.912 ;
        RECT 0.6 0.648 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
      LAYER V0 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.324 0.684 1.332 0.756 ;
        RECT 0.324 0.252 0.544 0.324 ;
        RECT 0.324 0.252 0.396 0.756 ;
      LAYER V0 ;
        RECT 0.324 0.612 0.396 0.684 ;
        RECT 0.396 0.252 0.468 0.324 ;
        RECT 1.26 0.684 1.332 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.108 0.684 0.18 ;
  END
END OAI211xp5_ASAP7_6t_fix

MACRO OAI21x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.372 1.224 0.608 ;
        RECT 0.58 0.684 1.152 0.756 ;
        RECT 1.08 0.536 1.152 0.756 ;
        RECT 0.428 0.252 0.66 0.324 ;
        RECT 0.58 0.536 0.652 0.756 ;
        RECT 0.504 0.536 0.652 0.608 ;
        RECT 0.504 0.252 0.576 0.608 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
        RECT 1.152 0.392 1.224 0.464 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.252 1.024 0.324 ;
        RECT 0.76 0.396 0.996 0.468 ;
        RECT 0.76 0.54 0.98 0.612 ;
        RECT 0.76 0.252 0.832 0.612 ;
      LAYER V0 ;
        RECT 0.924 0.396 0.996 0.468 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.288 0.396 1.44 0.468 ;
      LAYER M1 ;
        RECT 1.368 0.376 1.44 0.58 ;
        RECT 0.288 0.38 0.36 0.584 ;
      LAYER V1 ;
        RECT 0.288 0.396 0.36 0.468 ;
        RECT 1.368 0.396 1.44 0.468 ;
      LAYER V0 ;
        RECT 0.288 0.4 0.36 0.472 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.368 0.684 1.564 0.756 ;
      LAYER M1 ;
        RECT 1.26 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.476 0.108 1.656 0.18 ;
        RECT 0.072 0.684 0.468 0.756 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V1 ;
        RECT 0.388 0.684 0.46 0.756 ;
        RECT 1.268 0.684 1.34 0.756 ;
      LAYER V0 ;
        RECT 0.18 0.108 0.252 0.18 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.332 0.18 ;
  END
END OAI21x1_ASAP7_6t_fix

MACRO OAI21xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.508 0.144 0.58 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.472 0.564 0.544 ;
        RECT 0.288 0.684 0.488 0.756 ;
        RECT 0.288 0.304 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.492 0.472 0.564 0.544 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.688 0.54 0.836 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.46 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.468 0.792 0.54 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.816 -0.048 0.912 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.396 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.612 0.684 0.684 0.756 ;
    END
  END Y
END OAI21xp33_ASAP7_6t_fix

MACRO OAI21xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.068 0.684 0.216 0.756 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.412 0.6 0.484 ;
        RECT 0.34 0.684 0.488 0.756 ;
        RECT 0.36 0.412 0.432 0.756 ;
      LAYER V0 ;
        RECT 0.508 0.412 0.58 0.484 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.868 0.608 1.016 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.86 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.684 0.792 0.756 ;
        RECT 0.72 0.252 0.792 0.756 ;
        RECT 0.364 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.384 0.252 0.456 0.324 ;
        RECT 0.612 0.684 0.684 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.108 0.684 0.18 ;
  END
END OAI21xp5_ASAP7_6t_fix

MACRO OAI221xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.396 1.484 0.468 ;
        RECT 1.152 0.54 1.372 0.612 ;
        RECT 1.152 0.396 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.468 1.224 0.54 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.108 1.872 0.728 ;
        RECT 1.692 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.396 0.62 0.468 ;
        RECT 0.072 0.54 0.292 0.612 ;
        RECT 0.072 0.396 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.216 0.396 0.288 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.416 0.54 0.82 0.612 ;
        RECT 0.748 0.424 0.82 0.612 ;
      LAYER V0 ;
        RECT 0.748 0.468 0.82 0.54 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 1.008 0.756 ;
        RECT 0.936 0.424 1.008 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.468 1.008 0.54 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.464 0.648 1.56 0.912 ;
        RECT 0.816 0.648 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.728 0.828 1.8 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.728 -0.036 1.8 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.656 0.756 ;
        RECT 1.584 0.252 1.656 0.756 ;
        RECT 0.072 0.252 1.656 0.324 ;
      LAYER V0 ;
        RECT 0.072 0.252 0.144 0.324 ;
        RECT 0.612 0.252 0.684 0.324 ;
        RECT 1.26 0.684 1.332 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.108 1.548 0.18 ;
      RECT 0.396 0.108 0.9 0.18 ;
  END
END OAI221xp5_ASAP7_6t_fix

MACRO OAI222xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222xp33_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.144 0.728 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.54 0.62 0.612 ;
        RECT 0.376 0.396 0.596 0.468 ;
        RECT 0.376 0.396 0.448 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.288 0.684 1.44 0.756 ;
        RECT 1.368 0.396 1.44 0.756 ;
        RECT 1.132 0.396 1.44 0.468 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.804 0.54 1.024 0.612 ;
        RECT 0.952 0.396 1.024 0.612 ;
        RECT 0.72 0.396 1.024 0.468 ;
      LAYER V0 ;
        RECT 0.74 0.396 0.812 0.468 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.684 1.816 0.756 ;
        RECT 1.584 0.252 1.732 0.324 ;
        RECT 1.584 0.252 1.656 0.756 ;
      LAYER V0 ;
        RECT 1.584 0.4 1.656 0.472 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.684 2.088 0.756 ;
        RECT 2.016 0.108 2.088 0.756 ;
        RECT 1.888 0.108 2.088 0.18 ;
      LAYER V0 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.224 0.684 1.14 0.756 ;
        RECT 0.224 0.252 0.452 0.324 ;
        RECT 0.224 0.252 0.296 0.756 ;
      LAYER V0 ;
        RECT 0.352 0.252 0.424 0.324 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 1.044 0.684 1.116 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.856 0.252 1.44 0.324 ;
      RECT 1.368 0.108 1.44 0.324 ;
      RECT 1.368 0.108 1.764 0.18 ;
      RECT 0.18 0.108 1.136 0.18 ;
  END
END OAI222xp33_ASAP7_6t_fix

MACRO OAI22x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.06 0.396 1.568 0.468 ;
      LAYER M1 ;
        RECT 1.44 0.396 1.588 0.468 ;
        RECT 0.068 0.252 0.216 0.612 ;
      LAYER V1 ;
        RECT 0.08 0.396 0.152 0.468 ;
        RECT 1.476 0.396 1.548 0.468 ;
      LAYER V0 ;
        RECT 1.476 0.396 1.548 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.732 0.408 1.896 0.48 ;
        RECT 1.124 0.54 1.804 0.612 ;
        RECT 1.732 0.408 1.804 0.612 ;
        RECT 1.124 0.408 1.196 0.612 ;
      LAYER V0 ;
        RECT 1.124 0.408 1.196 0.48 ;
        RECT 1.804 0.408 1.876 0.48 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.68 0.252 0.86 0.324 ;
        RECT 0.572 0.396 0.752 0.468 ;
        RECT 0.68 0.252 0.752 0.468 ;
      LAYER V0 ;
        RECT 0.608 0.396 0.68 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.54 1.008 0.612 ;
        RECT 0.936 0.4 1.008 0.612 ;
        RECT 0.288 0.252 0.468 0.324 ;
        RECT 0.288 0.252 0.36 0.612 ;
      LAYER V0 ;
        RECT 0.288 0.4 0.36 0.472 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.152 0.684 2.088 0.756 ;
        RECT 2.016 0.252 2.088 0.756 ;
        RECT 1.272 0.252 2.088 0.324 ;
      LAYER V0 ;
        RECT 0.18 0.684 0.252 0.756 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.292 0.252 1.364 0.324 ;
        RECT 1.66 0.252 1.732 0.324 ;
        RECT 1.908 0.684 1.98 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 2 0.18 ;
  END
END OAI22x1_ASAP7_6t_fix

MACRO OAI22xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.508 0.576 0.58 ;
        RECT 0.216 0.508 0.504 0.612 ;
        RECT 0.216 0.252 0.48 0.324 ;
        RECT 0.216 0.252 0.288 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.508 0.576 0.58 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.108 1.032 0.18 ;
        RECT 0.7 0.504 0.864 0.576 ;
        RECT 0.792 0.108 0.864 0.576 ;
      LAYER V0 ;
        RECT 0.72 0.504 0.792 0.576 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.684 1.44 0.756 ;
        RECT 1.368 0.108 1.44 0.756 ;
        RECT 1.22 0.108 1.44 0.18 ;
        RECT 1.152 0.488 1.224 0.756 ;
      LAYER V0 ;
        RECT 1.152 0.508 1.224 0.58 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.224 0.324 ;
        RECT 0.86 0.684 1.008 0.756 ;
        RECT 0.936 0.252 1.008 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.488 1.008 0.56 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.032 -0.048 1.128 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.684 0.756 ;
        RECT 0.072 0.108 0.684 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 0.612 0.108 0.684 0.18 ;
    END
  END Y
END OAI22xp33_ASAP7_6t_fix

MACRO OAI22xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.356 0.684 0.576 0.756 ;
        RECT 0.504 0.252 0.576 0.756 ;
        RECT 0.356 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.656 0.756 ;
        RECT 1.584 0.252 1.656 0.756 ;
        RECT 1.508 0.252 1.656 0.324 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.54 1.444 0.612 ;
        RECT 1.152 0.252 1.384 0.324 ;
        RECT 1.152 0.252 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.4 1.224 0.472 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.756 0.684 1.116 0.756 ;
        RECT 0.756 0.252 0.92 0.324 ;
        RECT 0.756 0.252 0.828 0.756 ;
      LAYER V0 ;
        RECT 0.828 0.252 0.9 0.324 ;
        RECT 1.044 0.684 1.116 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.108 1.548 0.18 ;
  END
END OAI22xp5_ASAP7_6t_fix

MACRO OAI311xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI311xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.68 0.54 0.828 0.612 ;
        RECT 0.68 0.252 0.828 0.324 ;
        RECT 0.72 0.252 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.684 0.576 0.756 ;
        RECT 0.504 0.252 0.576 0.756 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.14 0.684 0.288 0.756 ;
        RECT 0.216 0.108 0.288 0.756 ;
        RECT 0.14 0.108 0.288 0.18 ;
      LAYER V0 ;
        RECT 0.216 0.396 0.288 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.54 1.084 0.612 ;
        RECT 0.936 0.252 1.084 0.324 ;
        RECT 0.936 0.252 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.22 0.108 1.292 0.488 ;
        RECT 1.144 0.108 1.292 0.18 ;
      LAYER V0 ;
        RECT 1.22 0.396 1.292 0.468 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.68 0.684 1.44 0.756 ;
        RECT 1.368 0.18 1.44 0.756 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.368 0.18 1.44 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 0.9 0.18 ;
  END
END OAI311xp33_ASAP7_6t_fix

MACRO OAI31xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.684 1.008 0.756 ;
        RECT 0.936 0.252 1.008 0.756 ;
        RECT 0.812 0.252 1.008 0.324 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.416 0.684 0.576 0.756 ;
        RECT 0.504 0.252 0.576 0.756 ;
        RECT 0.372 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.292 0.756 ;
        RECT 0.072 0.112 0.22 0.184 ;
        RECT 0.072 0.112 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.484 0.324 ;
        RECT 1.152 0.54 1.3 0.612 ;
        RECT 1.152 0.252 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.648 1.56 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.396 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.372 0.108 0.9 0.18 ;
  END
END OAI31xp33_ASAP7_6t_fix

MACRO OAI321xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI321xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.676 0.252 0.824 0.324 ;
        RECT 0.72 0.252 0.792 0.472 ;
      LAYER V0 ;
        RECT 0.72 0.4 0.792 0.472 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.684 0.576 0.756 ;
        RECT 0.504 0.252 0.576 0.756 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.4 0.576 0.472 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.112 0.22 0.184 ;
        RECT 0.072 0.112 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.108 0.54 1.256 0.612 ;
        RECT 1.152 0.448 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.468 1.224 0.54 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.54 1.66 0.612 ;
        RECT 1.512 0.252 1.66 0.324 ;
        RECT 1.512 0.252 1.584 0.612 ;
      LAYER V0 ;
        RECT 1.512 0.396 1.584 0.468 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.136 0.324 ;
        RECT 0.86 0.54 1.008 0.612 ;
        RECT 0.936 0.252 1.008 0.612 ;
      LAYER V0 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.032 0.648 1.128 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 1.596 0.756 ;
        RECT 1.368 0.252 1.44 0.756 ;
        RECT 1.26 0.252 1.44 0.324 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 1.26 0.252 1.332 0.324 ;
        RECT 1.476 0.684 1.548 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.108 1.548 0.18 ;
      RECT 0.396 0.108 0.9 0.18 ;
  END
END OAI321xp33_ASAP7_6t_fix

MACRO OAI322xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI322xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.868 0.452 1.012 0.524 ;
        RECT 0.792 0.684 0.94 0.756 ;
        RECT 0.868 0.452 0.94 0.756 ;
      LAYER V0 ;
        RECT 0.94 0.452 1.012 0.524 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.168 0.252 1.316 0.324 ;
        RECT 1.136 0.54 1.284 0.612 ;
        RECT 1.168 0.252 1.24 0.612 ;
      LAYER V0 ;
        RECT 1.168 0.408 1.24 0.48 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.684 0.548 0.756 ;
        RECT 0.476 0.388 0.548 0.756 ;
        RECT 0.216 0.46 0.288 0.756 ;
      LAYER V0 ;
        RECT 0.476 0.408 0.548 0.48 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.684 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.264 1.872 0.728 ;
      LAYER V0 ;
        RECT 1.8 0.396 1.872 0.468 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 1.728 0.756 ;
        RECT 1.656 0.252 1.728 0.756 ;
        RECT 1.504 0.252 1.728 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.524 0.252 1.596 0.324 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.496 0.396 0.74 0.468 ;
      LAYER M1 ;
        RECT 0.62 0.396 0.768 0.468 ;
        RECT 0.62 0.396 0.692 0.684 ;
      LAYER V1 ;
        RECT 0.648 0.396 0.72 0.468 ;
      LAYER V0 ;
        RECT 0.696 0.396 0.768 0.468 ;
    END
  END A1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.416 0.396 1.66 0.468 ;
      LAYER M1 ;
        RECT 1.364 0.396 1.556 0.468 ;
      LAYER V1 ;
        RECT 1.436 0.396 1.508 0.468 ;
      LAYER V0 ;
        RECT 1.364 0.396 1.436 0.468 ;
    END
  END C2
  OBS
    LAYER M1 ;
      RECT 0.6 0.252 1.068 0.324 ;
      RECT 0.6 0.108 0.672 0.324 ;
      RECT 0.072 0.108 0.672 0.18 ;
      RECT 0.808 0.108 1.764 0.18 ;
  END
END OAI322xp33_ASAP7_6t_fix

MACRO OAI32xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.32 0.396 0.596 0.468 ;
        RECT 0.32 0.252 0.54 0.324 ;
        RECT 0.32 0.684 0.468 0.756 ;
        RECT 0.32 0.252 0.392 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.728 0.54 0.928 0.612 ;
        RECT 0.856 0.252 0.928 0.612 ;
        RECT 0.728 0.252 0.928 0.324 ;
      LAYER V0 ;
        RECT 0.856 0.396 0.928 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.028 0.54 1.296 0.612 ;
        RECT 1.224 0.252 1.296 0.612 ;
        RECT 1.028 0.252 1.296 0.324 ;
      LAYER V0 ;
        RECT 1.224 0.396 1.296 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.42 0.396 1.7 0.468 ;
        RECT 1.42 0.54 1.64 0.612 ;
        RECT 1.42 0.396 1.492 0.612 ;
      LAYER V0 ;
        RECT 1.608 0.396 1.68 0.468 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 0.816 0.54 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.684 1.872 0.756 ;
        RECT 1.8 0.252 1.872 0.756 ;
        RECT 1.456 0.252 1.872 0.324 ;
      LAYER V0 ;
        RECT 0.612 0.684 0.684 0.756 ;
        RECT 1.476 0.252 1.548 0.324 ;
        RECT 1.692 0.684 1.764 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.764 0.18 ;
  END
END OAI32xp33_ASAP7_6t_fix

MACRO OAI331xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI331xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.616 0.684 0.764 0.756 ;
        RECT 0.692 0.388 0.764 0.756 ;
      LAYER V0 ;
        RECT 0.692 0.408 0.764 0.48 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.444 0.576 0.516 ;
        RECT 0.356 0.684 0.504 0.756 ;
        RECT 0.432 0.252 0.504 0.756 ;
        RECT 0.356 0.252 0.504 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.444 0.576 0.516 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.836 0.684 1.008 0.756 ;
        RECT 0.836 0.396 0.984 0.468 ;
        RECT 0.836 0.396 0.908 0.756 ;
      LAYER V0 ;
        RECT 0.912 0.396 0.984 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.176 0.396 1.324 0.612 ;
        RECT 1.104 0.516 1.324 0.588 ;
      LAYER V0 ;
        RECT 1.104 0.516 1.176 0.588 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.396 0.54 1.664 0.612 ;
        RECT 1.396 0.388 1.468 0.612 ;
      LAYER V0 ;
        RECT 1.396 0.408 1.468 0.48 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.62 0.396 1.872 0.468 ;
        RECT 1.8 0.108 1.872 0.468 ;
        RECT 1.696 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.62 0.396 1.692 0.468 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.872 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.848 0.252 1.348 0.324 ;
      RECT 0.848 0.108 0.92 0.324 ;
      RECT 0.396 0.108 0.92 0.18 ;
      RECT 1.044 0.108 1.548 0.18 ;
  END
END OAI331xp33_ASAP7_6t_fix

MACRO OAI332xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI332xp33_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.692 0.252 0.764 0.56 ;
        RECT 0.6 0.252 0.764 0.324 ;
      LAYER V0 ;
        RECT 0.692 0.408 0.764 0.48 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.684 0.576 0.756 ;
        RECT 0.504 0.44 0.576 0.756 ;
        RECT 0.288 0.252 0.452 0.324 ;
        RECT 0.288 0.252 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.44 0.576 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.468 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.836 0.408 0.984 0.48 ;
        RECT 0.744 0.684 0.908 0.756 ;
        RECT 0.836 0.388 0.908 0.756 ;
      LAYER V0 ;
        RECT 0.912 0.408 0.984 0.48 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.084 0.444 1.232 0.516 ;
        RECT 1.008 0.684 1.156 0.756 ;
        RECT 1.084 0.444 1.156 0.756 ;
      LAYER V0 ;
        RECT 1.16 0.444 1.232 0.516 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.252 2.088 0.728 ;
      LAYER V0 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.684 1.944 0.756 ;
        RECT 1.872 0.252 1.944 0.756 ;
        RECT 1.72 0.252 1.944 0.324 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.74 0.252 1.812 0.324 ;
    END
  END Y
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.36 0.396 1.668 0.468 ;
      LAYER M1 ;
        RECT 1.432 0.396 1.504 0.584 ;
        RECT 1.356 0.396 1.504 0.468 ;
      LAYER V1 ;
        RECT 1.396 0.396 1.468 0.468 ;
      LAYER V0 ;
        RECT 1.356 0.396 1.428 0.468 ;
    END
  END B3
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.44 0.54 1.736 0.612 ;
      LAYER M1 ;
        RECT 1.576 0.54 1.724 0.612 ;
        RECT 1.576 0.408 1.648 0.612 ;
      LAYER V1 ;
        RECT 1.636 0.54 1.708 0.612 ;
      LAYER V0 ;
        RECT 1.576 0.408 1.648 0.48 ;
    END
  END C2
  OBS
    LAYER M1 ;
      RECT 1.024 0.252 1.548 0.324 ;
      RECT 1.476 0.108 1.548 0.324 ;
      RECT 1.476 0.108 1.98 0.18 ;
      RECT 0.396 0.108 1.332 0.18 ;
  END
END OAI332xp33_ASAP7_6t_fix

MACRO OAI333xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI333xp33_ASAP7_6t_fix 0 0 ;
  SIZE 2.808 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.592 0.684 2.74 0.756 ;
        RECT 2.592 0.396 2.74 0.468 ;
        RECT 2.592 0.396 2.664 0.756 ;
      LAYER V0 ;
        RECT 2.668 0.396 2.74 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.856 0.54 2.332 0.612 ;
        RECT 2.26 0.424 2.332 0.612 ;
      LAYER V0 ;
        RECT 2.26 0.444 2.332 0.516 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.836 0.396 2.068 0.468 ;
        RECT 1.836 0.252 2.056 0.324 ;
        RECT 1.836 0.252 1.908 0.468 ;
      LAYER V0 ;
        RECT 1.996 0.396 2.068 0.468 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.864 0.396 1.052 0.468 ;
        RECT 0.504 0.684 0.936 0.756 ;
        RECT 0.864 0.396 0.936 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.396 1.484 0.468 ;
        RECT 1.152 0.54 1.372 0.612 ;
        RECT 1.152 0.396 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.252 1.736 0.324 ;
        RECT 1.584 0.54 1.732 0.612 ;
        RECT 1.584 0.252 1.656 0.612 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.244 0.54 0.764 0.612 ;
        RECT 0.692 0.396 0.764 0.612 ;
      LAYER V0 ;
        RECT 0.692 0.396 0.764 0.468 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.396 0.548 0.468 ;
        RECT 0.216 0.252 0.436 0.324 ;
        RECT 0.216 0.252 0.288 0.468 ;
      LAYER V0 ;
        RECT 0.476 0.396 0.548 0.468 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.38 0.756 ;
        RECT 0.072 0.136 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.808 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.808 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.808 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.18 0.252 2.74 0.324 ;
        RECT 1.044 0.684 2.52 0.756 ;
        RECT 2.448 0.252 2.52 0.756 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 2.18 0.252 2.252 0.324 ;
        RECT 2.34 0.684 2.412 0.756 ;
        RECT 2.668 0.252 2.74 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.252 1.44 0.324 ;
      RECT 0.828 0.108 0.9 0.324 ;
      RECT 0.396 0.108 0.9 0.18 ;
      RECT 2.34 0.108 2.488 0.18 ;
      RECT 1.044 0.108 1.98 0.18 ;
    LAYER M2 ;
      RECT 1.9 0.108 2.452 0.18 ;
    LAYER V1 ;
      RECT 2.36 0.108 2.432 0.18 ;
      RECT 1.9 0.108 1.972 0.18 ;
  END
END OAI333xp33_ASAP7_6t_fix

MACRO OAI33xp33_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33xp33_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.504 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.504 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.684 1.304 0.756 ;
        RECT 1.152 0.284 1.304 0.356 ;
        RECT 1.152 0.284 1.224 0.756 ;
      LAYER V0 ;
        RECT 1.152 0.372 1.224 0.444 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.896 0.684 1.08 0.756 ;
        RECT 1.008 0.284 1.08 0.756 ;
        RECT 0.896 0.284 1.08 0.356 ;
      LAYER V0 ;
        RECT 0.936 0.284 1.008 0.356 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.608 0.216 0.756 ;
        RECT 0.072 0.396 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.576 0.684 0.748 0.756 ;
        RECT 0.576 0.408 0.648 0.756 ;
        RECT 0.484 0.408 0.648 0.48 ;
      LAYER V0 ;
        RECT 0.504 0.408 0.576 0.48 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.216 ;
        RECT 1.032 -0.048 1.128 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.252 0.648 0.324 ;
        RECT 0.288 0.684 0.468 0.756 ;
        RECT 0.288 0.252 0.36 0.756 ;
        RECT 0.18 0.18 0.252 0.324 ;
      LAYER V0 ;
        RECT 0.18 0.18 0.252 0.252 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.576 0.252 0.648 0.324 ;
    END
  END Y
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.728 0.396 1.448 0.468 ;
      LAYER M1 ;
        RECT 0.748 0.5 0.896 0.572 ;
        RECT 0.748 0.388 0.82 0.572 ;
      LAYER V1 ;
        RECT 0.748 0.396 0.82 0.468 ;
      LAYER V0 ;
        RECT 0.748 0.408 0.82 0.48 ;
    END
  END B3
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.332 0.18 ;
  END
END OAI33xp33_ASAP7_6t_fix

MACRO OR2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.28 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.28 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.08 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.08 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.08 0.048 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 1.008 0.756 ;
        RECT 0.936 0.108 1.008 0.756 ;
        RECT 0.828 0.108 1.008 0.18 ;
      LAYER V0 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.72 0.756 ;
      RECT 0.648 0.108 0.72 0.756 ;
      RECT 0.648 0.396 0.836 0.468 ;
      RECT 0.396 0.108 0.72 0.18 ;
  END
END OR2x1_ASAP7_6t_fix

MACRO OR2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.584 ;
        RECT 0.288 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.36 0.612 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 0.828 0.108 1.224 0.18 ;
        RECT 0.828 0.592 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.272 ;
      LAYER V0 ;
        RECT 0.828 0.612 0.9 0.684 ;
        RECT 0.828 0.18 0.9 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.684 0.72 0.756 ;
      RECT 0.648 0.108 0.72 0.756 ;
      RECT 0.648 0.396 0.812 0.468 ;
      RECT 0.396 0.108 0.72 0.18 ;
  END
END OR2x2_ASAP7_6t_fix

MACRO OR2x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x4_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.352 0.54 0.576 0.612 ;
        RECT 0.504 0.252 0.576 0.612 ;
        RECT 0.352 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.224 0.756 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.684 1.584 0.756 ;
        RECT 1.512 0.108 1.584 0.756 ;
        RECT 0.828 0.108 1.584 0.18 ;
        RECT 1.26 0.592 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.272 ;
        RECT 0.828 0.592 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.272 ;
      LAYER V0 ;
        RECT 0.828 0.612 0.9 0.684 ;
        RECT 0.828 0.18 0.9 0.252 ;
        RECT 1.26 0.612 1.332 0.684 ;
        RECT 1.26 0.18 1.332 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.684 0.72 0.756 ;
      RECT 0.648 0.108 0.72 0.756 ;
      RECT 0.648 0.396 0.812 0.468 ;
      RECT 0.376 0.108 0.72 0.18 ;
  END
END OR2x4_ASAP7_6t_fix

MACRO OR2x6_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x6_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.324 0.576 0.396 ;
        RECT 0.288 0.54 0.504 0.612 ;
        RECT 0.432 0.324 0.504 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.324 0.576 0.396 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 1.008 0.756 ;
        RECT 0.936 0.376 1.008 0.756 ;
        RECT 0.072 0.108 0.224 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.328 0.54 2.424 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.328 -0.048 2.424 0.324 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.684 2.216 0.756 ;
        RECT 1.24 0.108 2.216 0.18 ;
        RECT 1.8 0.108 1.872 0.756 ;
      LAYER V0 ;
        RECT 1.26 0.684 1.332 0.756 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 2.124 0.684 2.196 0.756 ;
        RECT 2.124 0.108 2.196 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.54 0.792 0.612 ;
      RECT 0.72 0.108 0.792 0.612 ;
      RECT 1.08 0.396 1.244 0.468 ;
      RECT 1.08 0.204 1.152 0.468 ;
      RECT 0.9 0.204 1.152 0.276 ;
      RECT 0.9 0.108 0.972 0.276 ;
      RECT 0.376 0.108 0.972 0.18 ;
  END
END OR2x6_ASAP7_6t_fix

MACRO OR3x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.224 0.756 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.38 0.576 0.452 ;
        RECT 0.356 0.684 0.504 0.756 ;
        RECT 0.432 0.28 0.504 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.38 0.576 0.452 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.616 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.644 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.296 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.296 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.296 0.048 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 1.224 0.756 ;
        RECT 1.152 0.108 1.224 0.756 ;
        RECT 1.044 0.108 1.224 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.044 0.108 1.116 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.864 0.396 1.028 0.468 ;
      RECT 0.156 0.108 0.936 0.18 ;
  END
END OR3x1_ASAP7_6t_fix

MACRO OR3x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.288 0.612 ;
        RECT 0.072 0.28 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.396 0.576 0.468 ;
        RECT 0.432 0.252 0.504 0.584 ;
        RECT 0.32 0.252 0.504 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.54 0.792 0.612 ;
        RECT 0.72 0.252 0.792 0.612 ;
        RECT 0.644 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.512 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.512 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.512 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.54 1.44 0.612 ;
        RECT 1.368 0.252 1.44 0.612 ;
        RECT 1.044 0.252 1.44 0.324 ;
        RECT 1.044 0.54 1.116 0.728 ;
        RECT 1.044 0.136 1.116 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.636 1.116 0.708 ;
        RECT 1.044 0.156 1.116 0.228 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.156 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.864 0.396 1.116 0.468 ;
      RECT 0.156 0.108 0.936 0.18 ;
  END
END OR3x2_ASAP7_6t_fix

MACRO OR3x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x4_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.296 0.612 ;
        RECT 0.072 0.252 0.296 0.324 ;
        RECT 0.072 0.252 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.42 0.576 0.492 ;
        RECT 0.28 0.684 0.504 0.756 ;
        RECT 0.432 0.28 0.504 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.42 0.576 0.492 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.792 0.536 ;
        RECT 0.64 0.252 0.792 0.324 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.816 0.54 0.912 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.324 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.54 1.872 0.612 ;
        RECT 1.8 0.232 1.872 0.612 ;
        RECT 1.044 0.252 1.872 0.324 ;
        RECT 1.476 0.232 1.872 0.324 ;
        RECT 1.476 0.54 1.548 0.728 ;
        RECT 1.476 0.136 1.548 0.324 ;
        RECT 1.044 0.54 1.116 0.728 ;
        RECT 1.044 0.136 1.116 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.636 1.116 0.708 ;
        RECT 1.044 0.156 1.116 0.228 ;
        RECT 1.476 0.636 1.548 0.708 ;
        RECT 1.476 0.156 1.548 0.228 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.684 0.936 0.756 ;
      RECT 0.864 0.108 0.936 0.756 ;
      RECT 0.864 0.396 1.228 0.468 ;
      RECT 0.156 0.108 0.936 0.18 ;
  END
END OR3x4_ASAP7_6t_fix

MACRO OR4x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.54 0.308 0.612 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.684 0.548 0.756 ;
        RECT 0.476 0.252 0.548 0.756 ;
        RECT 0.4 0.252 0.548 0.324 ;
      LAYER V0 ;
        RECT 0.476 0.396 0.548 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.54 0.864 0.612 ;
        RECT 0.644 0.396 0.864 0.468 ;
        RECT 0.644 0.252 0.864 0.324 ;
        RECT 0.644 0.252 0.716 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.964 0.54 1.184 0.612 ;
        RECT 0.964 0.252 1.184 0.324 ;
        RECT 0.964 0.252 1.036 0.612 ;
      LAYER V0 ;
        RECT 0.964 0.396 1.036 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.684 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.456 0.108 1.656 0.18 ;
      LAYER V0 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.476 0.108 1.548 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.684 1.356 0.756 ;
      RECT 1.284 0.108 1.356 0.756 ;
      RECT 0.396 0.108 1.356 0.18 ;
  END
END OR4x1_ASAP7_6t_fix

MACRO OR4x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.064 0.536 0.288 0.608 ;
        RECT 0.216 0.108 0.288 0.608 ;
        RECT 0.064 0.108 0.288 0.18 ;
      LAYER V0 ;
        RECT 0.216 0.396 0.288 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.684 0.576 0.756 ;
        RECT 0.504 0.28 0.576 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.54 0.868 0.612 ;
        RECT 0.648 0.464 0.792 0.612 ;
        RECT 0.72 0.392 0.792 0.612 ;
      LAYER V0 ;
        RECT 0.72 0.392 0.792 0.464 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.488 ;
        RECT 0.86 0.252 1.008 0.324 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.54 1.656 0.612 ;
        RECT 1.584 0.252 1.656 0.612 ;
        RECT 1.26 0.252 1.656 0.324 ;
        RECT 1.26 0.54 1.332 0.728 ;
        RECT 1.26 0.136 1.332 0.324 ;
      LAYER V0 ;
        RECT 1.26 0.636 1.332 0.708 ;
        RECT 1.26 0.156 1.332 0.228 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.684 1.152 0.756 ;
      RECT 1.08 0.108 1.152 0.756 ;
      RECT 1.08 0.396 1.344 0.468 ;
      RECT 0.396 0.108 1.152 0.18 ;
  END
END OR4x2_ASAP7_6t_fix

MACRO OR4x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4x4_ASAP7_6t_fix 0 0 ;
  SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.252 1.872 0.584 ;
        RECT 1.576 0.252 1.872 0.324 ;
      LAYER V0 ;
        RECT 1.8 0.388 1.872 0.46 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.684 1.784 0.756 ;
        RECT 1.584 0.444 1.656 0.756 ;
      LAYER V0 ;
        RECT 1.584 0.444 1.656 0.516 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.324 0.608 1.472 0.756 ;
        RECT 1.368 0.252 1.44 0.756 ;
        RECT 1.24 0.252 1.44 0.324 ;
      LAYER V0 ;
        RECT 1.368 0.388 1.44 0.46 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.02 0.404 1.224 0.476 ;
        RECT 1.02 0.608 1.168 0.756 ;
        RECT 1.02 0.404 1.092 0.756 ;
      LAYER V0 ;
        RECT 1.152 0.404 1.224 0.476 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.16 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.16 0.912 ;
        RECT 1.032 0.54 1.128 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.16 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 1.032 -0.048 1.128 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.684 0.92 0.756 ;
        RECT 0.288 0.108 0.9 0.18 ;
        RECT 0.288 0.108 0.36 0.756 ;
      LAYER V0 ;
        RECT 0.396 0.684 0.468 0.756 ;
        RECT 0.396 0.108 0.468 0.18 ;
        RECT 0.828 0.684 0.9 0.756 ;
        RECT 0.828 0.108 0.9 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.908 0.684 2.088 0.756 ;
      RECT 2.016 0.108 2.088 0.756 ;
      RECT 0.72 0.252 0.792 0.516 ;
      RECT 0.72 0.252 1.116 0.324 ;
      RECT 1.044 0.108 1.116 0.324 ;
      RECT 1.044 0.108 2.088 0.18 ;
  END
END OR4x4_ASAP7_6t_fix

MACRO OR5x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x1_ASAP7_6t_fix 0 0 ;
  SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.26 0.756 ;
        RECT 0.072 0.28 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.488 ;
        RECT 0.284 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.492 0.684 0.792 0.756 ;
        RECT 0.72 0.44 0.792 0.756 ;
      LAYER V0 ;
        RECT 0.72 0.44 0.792 0.512 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.488 ;
        RECT 0.82 0.252 1.008 0.324 ;
      LAYER V0 ;
        RECT 0.936 0.396 1.008 0.468 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.54 1.224 0.612 ;
        RECT 1.152 0.28 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.728 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.728 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.728 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.508 0.608 1.656 0.756 ;
        RECT 1.584 0.108 1.656 0.756 ;
        RECT 1.508 0.108 1.656 0.256 ;
      LAYER V0 ;
        RECT 1.584 0.396 1.656 0.468 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.684 1.432 0.756 ;
      RECT 1.36 0.108 1.432 0.756 ;
      RECT 0.16 0.108 1.432 0.18 ;
  END
END OR5x1_ASAP7_6t_fix

MACRO OR5x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x2_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.684 0.348 0.756 ;
        RECT 0.072 0.28 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.448 ;
        RECT 0.284 0.252 0.576 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.376 0.576 0.448 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5 0.684 0.792 0.756 ;
        RECT 0.72 0.396 0.792 0.756 ;
      LAYER V0 ;
        RECT 0.72 0.396 0.792 0.468 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.896 0.252 1.044 0.4 ;
        RECT 0.936 0.252 1.008 0.472 ;
      LAYER V0 ;
        RECT 0.936 0.4 1.008 0.472 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.244 0.54 1.18 0.612 ;
      LAYER M1 ;
        RECT 1.076 0.54 1.224 0.612 ;
        RECT 1.152 0.332 1.224 0.612 ;
        RECT 0.244 0.396 0.392 0.612 ;
      LAYER V1 ;
        RECT 0.288 0.54 0.36 0.612 ;
        RECT 1.088 0.54 1.16 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.396 1.224 0.468 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.684 1.736 0.756 ;
        RECT 1.512 0.108 1.736 0.18 ;
        RECT 1.512 0.108 1.584 0.756 ;
      LAYER V0 ;
        RECT 1.512 0.612 1.584 0.684 ;
        RECT 1.512 0.18 1.584 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.684 1.44 0.756 ;
      RECT 1.368 0.108 1.44 0.756 ;
      RECT 0.16 0.108 1.44 0.18 ;
  END
END OR5x2_ASAP7_6t_fix

MACRO OR5x4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5x4_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.684 0.36 0.756 ;
        RECT 0.288 0.252 0.36 0.756 ;
        RECT 0.068 0.252 0.36 0.324 ;
      LAYER V0 ;
        RECT 0.288 0.324 0.36 0.396 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.684 0.836 0.756 ;
        RECT 0.464 0.252 0.612 0.324 ;
        RECT 0.504 0.252 0.576 0.756 ;
      LAYER V0 ;
        RECT 0.504 0.444 0.576 0.516 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 1.052 0.324 ;
        RECT 0.72 0.252 0.792 0.584 ;
      LAYER V0 ;
        RECT 0.72 0.324 0.792 0.396 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.684 1.352 0.756 ;
        RECT 0.936 0.424 1.008 0.756 ;
      LAYER V0 ;
        RECT 0.936 0.444 1.008 0.516 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.54 2.096 0.612 ;
        RECT 1.152 0.28 1.224 0.612 ;
      LAYER V0 ;
        RECT 1.152 0.404 1.224 0.476 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.816 -0.048 0.912 0.216 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.684 2.304 0.756 ;
        RECT 2.232 0.108 2.304 0.756 ;
        RECT 1.476 0.108 2.304 0.18 ;
        RECT 1.476 0.108 1.548 0.296 ;
      LAYER V0 ;
        RECT 1.476 0.684 1.548 0.756 ;
        RECT 1.476 0.18 1.548 0.252 ;
        RECT 1.908 0.684 1.98 0.756 ;
        RECT 1.908 0.108 1.98 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.332 0.396 1.66 0.468 ;
      RECT 1.332 0.108 1.404 0.468 ;
      RECT 0.18 0.108 1.404 0.18 ;
  END
END OR5x4_ASAP7_6t_fix

MACRO SDFLx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx1_ASAP7_6t_fix 0 0 ;
  SIZE 6.048 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.684 0.396 0.756 ;
        RECT 0.324 0.252 0.396 0.756 ;
        RECT 0.068 0.252 0.396 0.324 ;
      LAYER V0 ;
        RECT 0.324 0.448 0.396 0.52 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.784 0.684 5.968 0.756 ;
        RECT 5.896 0.244 5.968 0.756 ;
      LAYER V0 ;
        RECT 5.896 0.564 5.968 0.636 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 6.048 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 6.048 0.912 ;
        RECT 5.568 0.54 5.664 0.912 ;
        RECT 4.488 0.648 4.584 0.912 ;
        RECT 3.408 0.648 3.504 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
        RECT 5.796 0.828 5.868 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.048 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 6.048 0.048 ;
        RECT 5.568 -0.048 5.664 0.324 ;
        RECT 4.488 -0.048 4.584 0.216 ;
        RECT 3.408 -0.048 3.504 0.216 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
        RECT 5.796 -0.036 5.868 0.036 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.028 0.54 2.94 0.612 ;
      LAYER M1 ;
        RECT 2.044 0.54 2.264 0.612 ;
        RECT 2.192 0.396 2.264 0.612 ;
        RECT 2.044 0.396 2.264 0.468 ;
      LAYER V1 ;
        RECT 2.052 0.54 2.124 0.612 ;
      LAYER V0 ;
        RECT 2.084 0.396 2.156 0.468 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.792 0.108 5.696 0.18 ;
      LAYER M1 ;
        RECT 5.596 0.108 5.816 0.18 ;
        RECT 5.472 0.38 5.668 0.452 ;
        RECT 5.596 0.108 5.668 0.452 ;
        RECT 0.936 0.108 1.008 0.276 ;
        RECT 0.808 0.108 1.008 0.18 ;
      LAYER V1 ;
        RECT 0.82 0.108 0.892 0.18 ;
        RECT 5.604 0.108 5.676 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.184 1.008 0.256 ;
        RECT 5.472 0.38 5.544 0.452 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.628 0.54 1.768 0.612 ;
      LAYER M1 ;
        RECT 1.656 0.54 1.804 0.612 ;
        RECT 1.656 0.38 1.728 0.612 ;
        RECT 1.364 0.38 1.728 0.452 ;
      LAYER V1 ;
        RECT 1.676 0.54 1.748 0.612 ;
      LAYER V0 ;
        RECT 1.58 0.38 1.656 0.452 ;
    END
  END SI
  OBS
    LAYER M1 ;
      RECT 5.364 0.684 5.6 0.756 ;
      RECT 5.528 0.54 5.6 0.756 ;
      RECT 5.38 0.54 5.608 0.612 ;
      RECT 4.048 0.684 4.8 0.756 ;
      RECT 4.728 0.108 4.8 0.756 ;
      RECT 5.264 0.108 5.336 0.332 ;
      RECT 4.048 0.108 5.336 0.18 ;
      RECT 4.14 0.54 4.656 0.612 ;
      RECT 4.584 0.252 4.656 0.612 ;
      RECT 4.14 0.468 4.212 0.612 ;
      RECT 4.436 0.252 4.656 0.324 ;
      RECT 3.792 0.52 3.992 0.592 ;
      RECT 3.92 0.272 3.992 0.592 ;
      RECT 3.92 0.272 4.232 0.344 ;
      RECT 2.988 0.684 3.528 0.756 ;
      RECT 3.456 0.108 3.528 0.756 ;
      RECT 2.752 0.108 3.528 0.18 ;
      RECT 3.22 0.54 3.368 0.612 ;
      RECT 3.296 0.28 3.368 0.612 ;
      RECT 2.88 0.252 2.952 0.468 ;
      RECT 2.804 0.252 2.952 0.324 ;
      RECT 2.74 0.608 2.888 0.756 ;
      RECT 2.336 0.54 2.812 0.612 ;
      RECT 2.336 0.252 2.408 0.612 ;
      RECT 1.824 0.252 1.896 0.456 ;
      RECT 1.824 0.252 2.408 0.324 ;
      RECT 0.976 0.54 1.124 0.756 ;
      RECT 0.976 0.54 1.5 0.612 ;
      RECT 0.504 0.108 0.576 0.364 ;
      RECT 0.156 0.108 0.576 0.18 ;
      RECT 5.74 0.288 5.812 0.476 ;
      RECT 4.98 0.308 5.052 0.496 ;
      RECT 4.336 0.396 4.484 0.468 ;
      RECT 3.76 0.136 3.832 0.352 ;
      RECT 3.616 0.144 3.688 0.72 ;
      RECT 3.096 0.288 3.168 0.476 ;
      RECT 2.608 0.396 2.756 0.468 ;
      RECT 2.34 0.684 2.492 0.756 ;
      RECT 1.24 0.108 2.216 0.18 ;
      RECT 1.26 0.684 2.216 0.756 ;
      RECT 0.688 0.36 0.76 0.508 ;
    LAYER M2 ;
      RECT 5.74 0.252 5.812 0.488 ;
      RECT 5.24 0.252 5.812 0.324 ;
      RECT 2.784 0.684 5.328 0.756 ;
      RECT 5.256 0.54 5.328 0.756 ;
      RECT 5.256 0.54 5.62 0.612 ;
      RECT 4.372 0.396 5.072 0.468 ;
      RECT 0.484 0.252 4.676 0.324 ;
      RECT 0.668 0.396 4.012 0.468 ;
      RECT 3.244 0.54 3.708 0.612 ;
      RECT 1.012 0.684 2.588 0.756 ;
    LAYER V1 ;
      RECT 5.74 0.396 5.812 0.468 ;
      RECT 5.528 0.54 5.6 0.612 ;
      RECT 5.264 0.252 5.336 0.324 ;
      RECT 4.98 0.396 5.052 0.468 ;
      RECT 4.576 0.252 4.648 0.324 ;
      RECT 4.392 0.396 4.464 0.468 ;
      RECT 3.92 0.396 3.992 0.468 ;
      RECT 3.76 0.252 3.832 0.324 ;
      RECT 3.616 0.54 3.688 0.612 ;
      RECT 3.264 0.54 3.336 0.612 ;
      RECT 3.096 0.396 3.168 0.468 ;
      RECT 2.816 0.252 2.888 0.324 ;
      RECT 2.804 0.684 2.876 0.756 ;
      RECT 2.676 0.396 2.748 0.468 ;
      RECT 2.388 0.684 2.46 0.756 ;
      RECT 1.04 0.684 1.112 0.756 ;
      RECT 0.688 0.396 0.76 0.468 ;
      RECT 0.504 0.252 0.576 0.324 ;
  END
END SDFLx1_ASAP7_6t_fix

MACRO SDFLx2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx2_ASAP7_6t_fix 0 0 ;
  SIZE 6.264 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.684 0.396 0.756 ;
        RECT 0.324 0.252 0.396 0.756 ;
        RECT 0.068 0.252 0.396 0.324 ;
      LAYER V0 ;
        RECT 0.324 0.448 0.396 0.52 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.828 0.54 2.148 0.612 ;
      LAYER M1 ;
        RECT 2.044 0.54 2.264 0.612 ;
        RECT 2.192 0.396 2.264 0.612 ;
        RECT 2.044 0.396 2.264 0.468 ;
      LAYER V1 ;
        RECT 2.052 0.54 2.124 0.612 ;
      LAYER V0 ;
        RECT 2.084 0.396 2.156 0.468 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.796 0.108 6 0.18 ;
        RECT 5.776 0.684 5.968 0.756 ;
        RECT 5.896 0.108 5.968 0.756 ;
      LAYER V0 ;
        RECT 5.796 0.684 5.868 0.756 ;
        RECT 5.796 0.108 5.868 0.18 ;
    END
  END QN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.54 1.804 0.612 ;
        RECT 1.656 0.38 1.728 0.612 ;
        RECT 0.832 0.38 1.728 0.452 ;
        RECT 0.504 0.684 0.904 0.756 ;
        RECT 0.832 0.38 0.904 0.756 ;
        RECT 0.504 0.488 0.576 0.756 ;
      LAYER V0 ;
        RECT 1.58 0.38 1.656 0.452 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 6.264 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 6.264 0.912 ;
        RECT 6 0.54 6.096 0.912 ;
        RECT 5.568 0.54 5.664 0.912 ;
        RECT 4.488 0.648 4.584 0.912 ;
        RECT 3.408 0.648 3.504 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
        RECT 5.796 0.828 5.868 0.9 ;
        RECT 6.012 0.828 6.084 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.264 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 6.264 0.048 ;
        RECT 6 -0.048 6.096 0.324 ;
        RECT 5.568 -0.048 5.664 0.324 ;
        RECT 4.488 -0.048 4.584 0.216 ;
        RECT 3.408 -0.048 3.504 0.216 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
        RECT 5.796 -0.036 5.868 0.036 ;
        RECT 6.012 -0.036 6.084 0.036 ;
    END
  END VSS
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.792 0.108 5.68 0.18 ;
      LAYER M1 ;
        RECT 5.472 0.38 5.668 0.452 ;
        RECT 5.596 0.108 5.668 0.452 ;
        RECT 5.464 0.108 5.668 0.18 ;
        RECT 0.936 0.108 1.008 0.276 ;
        RECT 0.808 0.108 1.008 0.18 ;
      LAYER V1 ;
        RECT 0.82 0.108 0.892 0.18 ;
        RECT 5.588 0.108 5.66 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.184 1.008 0.256 ;
        RECT 5.472 0.38 5.544 0.452 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 5.364 0.684 5.6 0.756 ;
      RECT 5.528 0.54 5.6 0.756 ;
      RECT 5.38 0.54 5.608 0.612 ;
      RECT 4.048 0.684 4.8 0.756 ;
      RECT 4.728 0.108 4.8 0.756 ;
      RECT 5.264 0.108 5.336 0.332 ;
      RECT 4.048 0.108 5.336 0.18 ;
      RECT 4.14 0.54 4.656 0.612 ;
      RECT 4.584 0.252 4.656 0.612 ;
      RECT 4.14 0.468 4.212 0.612 ;
      RECT 4.436 0.252 4.656 0.324 ;
      RECT 3.792 0.52 3.992 0.592 ;
      RECT 3.92 0.272 3.992 0.592 ;
      RECT 3.92 0.272 4.232 0.344 ;
      RECT 2.988 0.684 3.528 0.756 ;
      RECT 3.456 0.108 3.528 0.756 ;
      RECT 2.752 0.108 3.528 0.18 ;
      RECT 3.22 0.54 3.368 0.612 ;
      RECT 3.296 0.28 3.368 0.612 ;
      RECT 2.88 0.252 2.952 0.468 ;
      RECT 2.804 0.252 2.952 0.324 ;
      RECT 2.74 0.608 2.888 0.756 ;
      RECT 2.336 0.54 2.812 0.612 ;
      RECT 2.336 0.252 2.408 0.612 ;
      RECT 1.824 0.252 1.896 0.456 ;
      RECT 1.824 0.252 2.408 0.324 ;
      RECT 0.976 0.54 1.124 0.756 ;
      RECT 0.976 0.54 1.5 0.612 ;
      RECT 0.504 0.108 0.576 0.364 ;
      RECT 0.156 0.108 0.576 0.18 ;
      RECT 5.74 0.308 5.812 0.496 ;
      RECT 4.98 0.336 5.052 0.524 ;
      RECT 4.336 0.396 4.484 0.468 ;
      RECT 3.76 0.136 3.832 0.352 ;
      RECT 3.616 0.144 3.688 0.72 ;
      RECT 3.096 0.288 3.168 0.476 ;
      RECT 2.608 0.396 2.756 0.468 ;
      RECT 2.34 0.684 2.492 0.756 ;
      RECT 1.24 0.108 2.216 0.18 ;
      RECT 1.26 0.684 2.216 0.756 ;
      RECT 0.688 0.36 0.76 0.508 ;
    LAYER M2 ;
      RECT 5.74 0.252 5.812 0.488 ;
      RECT 5.24 0.252 5.812 0.324 ;
      RECT 2.784 0.684 5.328 0.756 ;
      RECT 5.256 0.54 5.328 0.756 ;
      RECT 5.256 0.54 5.62 0.612 ;
      RECT 4.372 0.396 5.072 0.468 ;
      RECT 0.484 0.252 4.676 0.324 ;
      RECT 0.668 0.396 4.012 0.468 ;
      RECT 3.244 0.54 3.708 0.612 ;
      RECT 1.012 0.684 2.588 0.756 ;
    LAYER V1 ;
      RECT 5.74 0.396 5.812 0.468 ;
      RECT 5.528 0.54 5.6 0.612 ;
      RECT 5.264 0.252 5.336 0.324 ;
      RECT 4.98 0.396 5.052 0.468 ;
      RECT 4.576 0.252 4.648 0.324 ;
      RECT 4.392 0.396 4.464 0.468 ;
      RECT 3.92 0.396 3.992 0.468 ;
      RECT 3.76 0.252 3.832 0.324 ;
      RECT 3.616 0.54 3.688 0.612 ;
      RECT 3.264 0.54 3.336 0.612 ;
      RECT 3.096 0.396 3.168 0.468 ;
      RECT 2.816 0.252 2.888 0.324 ;
      RECT 2.804 0.684 2.876 0.756 ;
      RECT 2.676 0.396 2.748 0.468 ;
      RECT 2.388 0.684 2.46 0.756 ;
      RECT 1.04 0.684 1.112 0.756 ;
      RECT 0.688 0.396 0.76 0.468 ;
      RECT 0.504 0.252 0.576 0.324 ;
  END
END SDFLx2_ASAP7_6t_fix

MACRO SDFLx3_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx3_ASAP7_6t_fix 0 0 ;
  SIZE 6.48 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.684 0.396 0.756 ;
        RECT 0.324 0.252 0.396 0.756 ;
        RECT 0.068 0.252 0.396 0.324 ;
      LAYER V0 ;
        RECT 0.324 0.448 0.396 0.52 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.828 0.54 2.148 0.612 ;
      LAYER M1 ;
        RECT 2.044 0.54 2.264 0.612 ;
        RECT 2.192 0.396 2.264 0.612 ;
        RECT 2.044 0.396 2.264 0.468 ;
      LAYER V1 ;
        RECT 2.052 0.54 2.124 0.612 ;
      LAYER V0 ;
        RECT 2.084 0.396 2.156 0.468 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.776 0.684 6.408 0.756 ;
        RECT 6.336 0.108 6.408 0.756 ;
        RECT 5.796 0.108 6.408 0.18 ;
      LAYER V0 ;
        RECT 5.796 0.684 5.868 0.756 ;
        RECT 5.796 0.108 5.868 0.18 ;
        RECT 6.228 0.684 6.3 0.756 ;
        RECT 6.228 0.108 6.3 0.18 ;
    END
  END QN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.54 1.804 0.612 ;
        RECT 1.656 0.38 1.728 0.612 ;
        RECT 0.832 0.38 1.728 0.452 ;
        RECT 0.504 0.684 0.904 0.756 ;
        RECT 0.832 0.38 0.904 0.756 ;
        RECT 0.504 0.488 0.576 0.756 ;
      LAYER V0 ;
        RECT 1.58 0.38 1.656 0.452 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 6.48 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 6.48 0.912 ;
        RECT 6 0.54 6.096 0.912 ;
        RECT 5.568 0.54 5.664 0.912 ;
        RECT 4.488 0.648 4.584 0.912 ;
        RECT 3.408 0.648 3.504 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
        RECT 5.796 0.828 5.868 0.9 ;
        RECT 6.012 0.828 6.084 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.48 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 6.48 0.048 ;
        RECT 6 -0.048 6.096 0.324 ;
        RECT 5.568 -0.048 5.664 0.324 ;
        RECT 4.488 -0.048 4.584 0.216 ;
        RECT 3.408 -0.048 3.504 0.216 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
        RECT 5.796 -0.036 5.868 0.036 ;
        RECT 6.012 -0.036 6.084 0.036 ;
    END
  END VSS
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.792 0.108 5.68 0.18 ;
      LAYER M1 ;
        RECT 5.472 0.38 5.668 0.452 ;
        RECT 5.596 0.108 5.668 0.452 ;
        RECT 5.464 0.108 5.668 0.18 ;
        RECT 0.936 0.108 1.008 0.276 ;
        RECT 0.808 0.108 1.008 0.18 ;
      LAYER V1 ;
        RECT 0.82 0.108 0.892 0.18 ;
        RECT 5.588 0.108 5.66 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.184 1.008 0.256 ;
        RECT 5.472 0.38 5.544 0.452 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 5.364 0.684 5.6 0.756 ;
      RECT 5.528 0.54 5.6 0.756 ;
      RECT 5.38 0.54 5.608 0.612 ;
      RECT 4.048 0.684 4.8 0.756 ;
      RECT 4.728 0.108 4.8 0.756 ;
      RECT 5.264 0.108 5.336 0.332 ;
      RECT 4.048 0.108 5.336 0.18 ;
      RECT 4.14 0.54 4.656 0.612 ;
      RECT 4.584 0.252 4.656 0.612 ;
      RECT 4.14 0.468 4.212 0.612 ;
      RECT 4.436 0.252 4.656 0.324 ;
      RECT 3.792 0.52 3.992 0.592 ;
      RECT 3.92 0.272 3.992 0.592 ;
      RECT 3.92 0.272 4.232 0.344 ;
      RECT 2.988 0.684 3.528 0.756 ;
      RECT 3.456 0.108 3.528 0.756 ;
      RECT 2.752 0.108 3.528 0.18 ;
      RECT 3.22 0.54 3.368 0.612 ;
      RECT 3.296 0.28 3.368 0.612 ;
      RECT 2.88 0.252 2.952 0.468 ;
      RECT 2.804 0.252 2.952 0.324 ;
      RECT 2.74 0.608 2.888 0.756 ;
      RECT 2.336 0.54 2.812 0.612 ;
      RECT 2.336 0.252 2.408 0.612 ;
      RECT 1.824 0.252 1.896 0.456 ;
      RECT 1.824 0.252 2.408 0.324 ;
      RECT 0.976 0.54 1.124 0.756 ;
      RECT 0.976 0.54 1.5 0.612 ;
      RECT 0.504 0.108 0.576 0.364 ;
      RECT 0.156 0.108 0.576 0.18 ;
      RECT 5.74 0.308 5.812 0.496 ;
      RECT 4.98 0.32 5.052 0.508 ;
      RECT 4.336 0.396 4.484 0.468 ;
      RECT 3.76 0.136 3.832 0.352 ;
      RECT 3.616 0.144 3.688 0.72 ;
      RECT 3.096 0.288 3.168 0.476 ;
      RECT 2.608 0.396 2.756 0.468 ;
      RECT 2.34 0.684 2.492 0.756 ;
      RECT 1.24 0.108 2.216 0.18 ;
      RECT 1.26 0.684 2.216 0.756 ;
      RECT 0.688 0.36 0.76 0.508 ;
    LAYER M2 ;
      RECT 5.74 0.252 5.812 0.488 ;
      RECT 5.24 0.252 5.812 0.324 ;
      RECT 2.784 0.684 5.328 0.756 ;
      RECT 5.256 0.54 5.328 0.756 ;
      RECT 5.256 0.54 5.62 0.612 ;
      RECT 4.372 0.396 5.072 0.468 ;
      RECT 0.484 0.252 4.676 0.324 ;
      RECT 0.668 0.396 4.012 0.468 ;
      RECT 3.244 0.54 3.708 0.612 ;
      RECT 1.012 0.684 2.588 0.756 ;
    LAYER V1 ;
      RECT 5.74 0.396 5.812 0.468 ;
      RECT 5.528 0.54 5.6 0.612 ;
      RECT 5.264 0.252 5.336 0.324 ;
      RECT 4.98 0.396 5.052 0.468 ;
      RECT 4.576 0.252 4.648 0.324 ;
      RECT 4.392 0.396 4.464 0.468 ;
      RECT 3.92 0.396 3.992 0.468 ;
      RECT 3.76 0.252 3.832 0.324 ;
      RECT 3.616 0.54 3.688 0.612 ;
      RECT 3.264 0.54 3.336 0.612 ;
      RECT 3.096 0.396 3.168 0.468 ;
      RECT 2.816 0.252 2.888 0.324 ;
      RECT 2.804 0.684 2.876 0.756 ;
      RECT 2.676 0.396 2.748 0.468 ;
      RECT 2.388 0.684 2.46 0.756 ;
      RECT 1.04 0.684 1.112 0.756 ;
      RECT 0.688 0.396 0.76 0.468 ;
      RECT 0.504 0.252 0.576 0.324 ;
  END
END SDFLx3_ASAP7_6t_fix

MACRO SDFLx4_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFLx4_ASAP7_6t_fix 0 0 ;
  SIZE 6.696 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.684 0.396 0.756 ;
        RECT 0.324 0.252 0.396 0.756 ;
        RECT 0.068 0.252 0.396 0.324 ;
      LAYER V0 ;
        RECT 0.324 0.448 0.396 0.52 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.828 0.54 2.148 0.612 ;
      LAYER M1 ;
        RECT 2.044 0.54 2.264 0.612 ;
        RECT 2.192 0.396 2.264 0.612 ;
        RECT 2.044 0.396 2.264 0.468 ;
      LAYER V1 ;
        RECT 2.052 0.54 2.124 0.612 ;
      LAYER V0 ;
        RECT 2.084 0.396 2.156 0.468 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.776 0.684 6.408 0.756 ;
        RECT 6.336 0.108 6.408 0.756 ;
        RECT 5.796 0.108 6.408 0.18 ;
      LAYER V0 ;
        RECT 5.796 0.684 5.868 0.756 ;
        RECT 5.796 0.108 5.868 0.18 ;
        RECT 6.228 0.684 6.3 0.756 ;
        RECT 6.228 0.108 6.3 0.18 ;
    END
  END QN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.54 1.804 0.612 ;
        RECT 1.656 0.38 1.728 0.612 ;
        RECT 0.832 0.38 1.728 0.452 ;
        RECT 0.504 0.684 0.904 0.756 ;
        RECT 0.832 0.38 0.904 0.756 ;
        RECT 0.504 0.488 0.576 0.756 ;
      LAYER V0 ;
        RECT 1.58 0.38 1.656 0.452 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 6.696 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 6.696 0.912 ;
        RECT 6.432 0.54 6.528 0.912 ;
        RECT 6 0.54 6.096 0.912 ;
        RECT 5.568 0.54 5.664 0.912 ;
        RECT 4.488 0.648 4.584 0.912 ;
        RECT 3.408 0.648 3.504 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
        RECT 2.556 0.828 2.628 0.9 ;
        RECT 2.772 0.828 2.844 0.9 ;
        RECT 2.988 0.828 3.06 0.9 ;
        RECT 3.204 0.828 3.276 0.9 ;
        RECT 3.42 0.828 3.492 0.9 ;
        RECT 3.636 0.828 3.708 0.9 ;
        RECT 3.852 0.828 3.924 0.9 ;
        RECT 4.068 0.828 4.14 0.9 ;
        RECT 4.284 0.828 4.356 0.9 ;
        RECT 4.5 0.828 4.572 0.9 ;
        RECT 4.716 0.828 4.788 0.9 ;
        RECT 4.932 0.828 5.004 0.9 ;
        RECT 5.148 0.828 5.22 0.9 ;
        RECT 5.364 0.828 5.436 0.9 ;
        RECT 5.58 0.828 5.652 0.9 ;
        RECT 5.796 0.828 5.868 0.9 ;
        RECT 6.012 0.828 6.084 0.9 ;
        RECT 6.228 0.828 6.3 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.696 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 6.696 0.048 ;
        RECT 6.432 -0.048 6.528 0.324 ;
        RECT 6 -0.048 6.096 0.324 ;
        RECT 5.568 -0.048 5.664 0.324 ;
        RECT 4.488 -0.048 4.584 0.216 ;
        RECT 3.408 -0.048 3.504 0.216 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
        RECT 2.556 -0.036 2.628 0.036 ;
        RECT 2.772 -0.036 2.844 0.036 ;
        RECT 2.988 -0.036 3.06 0.036 ;
        RECT 3.204 -0.036 3.276 0.036 ;
        RECT 3.42 -0.036 3.492 0.036 ;
        RECT 3.636 -0.036 3.708 0.036 ;
        RECT 3.852 -0.036 3.924 0.036 ;
        RECT 4.068 -0.036 4.14 0.036 ;
        RECT 4.284 -0.036 4.356 0.036 ;
        RECT 4.5 -0.036 4.572 0.036 ;
        RECT 4.716 -0.036 4.788 0.036 ;
        RECT 4.932 -0.036 5.004 0.036 ;
        RECT 5.148 -0.036 5.22 0.036 ;
        RECT 5.364 -0.036 5.436 0.036 ;
        RECT 5.58 -0.036 5.652 0.036 ;
        RECT 5.796 -0.036 5.868 0.036 ;
        RECT 6.012 -0.036 6.084 0.036 ;
        RECT 6.228 -0.036 6.3 0.036 ;
    END
  END VSS
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.792 0.108 5.68 0.18 ;
      LAYER M1 ;
        RECT 5.472 0.38 5.668 0.452 ;
        RECT 5.596 0.108 5.668 0.452 ;
        RECT 5.464 0.108 5.668 0.18 ;
        RECT 0.936 0.108 1.008 0.276 ;
        RECT 0.808 0.108 1.008 0.18 ;
      LAYER V1 ;
        RECT 0.82 0.108 0.892 0.18 ;
        RECT 5.588 0.108 5.66 0.18 ;
      LAYER V0 ;
        RECT 0.936 0.184 1.008 0.256 ;
        RECT 5.472 0.38 5.544 0.452 ;
    END
  END SE
  OBS
    LAYER M1 ;
      RECT 5.364 0.684 5.6 0.756 ;
      RECT 5.528 0.54 5.6 0.756 ;
      RECT 5.38 0.54 5.608 0.612 ;
      RECT 4.048 0.684 4.8 0.756 ;
      RECT 4.728 0.108 4.8 0.756 ;
      RECT 5.264 0.108 5.336 0.332 ;
      RECT 4.048 0.108 5.336 0.18 ;
      RECT 4.14 0.54 4.656 0.612 ;
      RECT 4.584 0.252 4.656 0.612 ;
      RECT 4.14 0.468 4.212 0.612 ;
      RECT 4.436 0.252 4.656 0.324 ;
      RECT 3.792 0.52 3.992 0.592 ;
      RECT 3.92 0.272 3.992 0.592 ;
      RECT 3.92 0.272 4.232 0.344 ;
      RECT 2.988 0.684 3.528 0.756 ;
      RECT 3.456 0.108 3.528 0.756 ;
      RECT 2.752 0.108 3.528 0.18 ;
      RECT 3.22 0.54 3.368 0.612 ;
      RECT 3.296 0.28 3.368 0.612 ;
      RECT 2.88 0.252 2.952 0.468 ;
      RECT 2.804 0.252 2.952 0.324 ;
      RECT 2.74 0.608 2.888 0.756 ;
      RECT 2.336 0.54 2.812 0.612 ;
      RECT 2.336 0.252 2.408 0.612 ;
      RECT 1.824 0.252 1.896 0.456 ;
      RECT 1.824 0.252 2.408 0.324 ;
      RECT 0.976 0.54 1.124 0.756 ;
      RECT 0.976 0.54 1.5 0.612 ;
      RECT 0.504 0.108 0.576 0.364 ;
      RECT 0.156 0.108 0.576 0.18 ;
      RECT 5.74 0.308 5.812 0.496 ;
      RECT 4.98 0.312 5.052 0.5 ;
      RECT 4.336 0.396 4.484 0.468 ;
      RECT 3.76 0.136 3.832 0.352 ;
      RECT 3.616 0.144 3.688 0.72 ;
      RECT 3.096 0.288 3.168 0.476 ;
      RECT 2.608 0.396 2.756 0.468 ;
      RECT 2.34 0.684 2.492 0.756 ;
      RECT 1.24 0.108 2.216 0.18 ;
      RECT 1.26 0.684 2.216 0.756 ;
      RECT 0.688 0.36 0.76 0.508 ;
    LAYER M2 ;
      RECT 5.74 0.252 5.812 0.488 ;
      RECT 5.24 0.252 5.812 0.324 ;
      RECT 2.784 0.684 5.328 0.756 ;
      RECT 5.256 0.54 5.328 0.756 ;
      RECT 5.256 0.54 5.62 0.612 ;
      RECT 4.372 0.396 5.072 0.468 ;
      RECT 0.484 0.252 4.676 0.324 ;
      RECT 0.668 0.396 4.012 0.468 ;
      RECT 3.244 0.54 3.708 0.612 ;
      RECT 1.012 0.684 2.588 0.756 ;
    LAYER V1 ;
      RECT 5.74 0.396 5.812 0.468 ;
      RECT 5.528 0.54 5.6 0.612 ;
      RECT 5.264 0.252 5.336 0.324 ;
      RECT 4.98 0.396 5.052 0.468 ;
      RECT 4.576 0.252 4.648 0.324 ;
      RECT 4.392 0.396 4.464 0.468 ;
      RECT 3.92 0.396 3.992 0.468 ;
      RECT 3.76 0.252 3.832 0.324 ;
      RECT 3.616 0.54 3.688 0.612 ;
      RECT 3.264 0.54 3.336 0.612 ;
      RECT 3.096 0.396 3.168 0.468 ;
      RECT 2.816 0.252 2.888 0.324 ;
      RECT 2.804 0.684 2.876 0.756 ;
      RECT 2.676 0.396 2.748 0.468 ;
      RECT 2.388 0.684 2.46 0.756 ;
      RECT 1.04 0.684 1.112 0.756 ;
      RECT 0.688 0.396 0.76 0.468 ;
      RECT 0.504 0.252 0.576 0.324 ;
  END
END SDFLx4_ASAP7_6t_fix

MACRO TAPCELL_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_ASAP7_6t_fix 0 0 ;
  SIZE 0.432 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.432 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.432 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.432 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.432 0.048 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
    END
  END VSS
END TAPCELL_ASAP7_6t_fix

MACRO TAPCELL_WITH_FILLER_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_WITH_FILLER_ASAP7_6t_fix 0 0 ;
  SIZE 0.648 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.648 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.648 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.648 0.048 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
    END
  END VSS
END TAPCELL_WITH_FILLER_ASAP7_6t_fix

MACRO TIEHIx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHIx1_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.324 0.684 0.576 0.756 ;
        RECT 0.504 0.272 0.576 0.756 ;
        RECT 0.268 0.272 0.576 0.344 ;
      LAYER V0 ;
        RECT 0.356 0.272 0.428 0.344 ;
        RECT 0.396 0.684 0.468 0.756 ;
    END
  END H
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.384 -0.048 0.48 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.072 0.52 0.336 0.592 ;
      RECT 0.072 0.108 0.144 0.592 ;
      RECT 0.072 0.108 0.324 0.18 ;
  END
END TIEHIx1_ASAP7_6t_fix

MACRO TIELOx1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELOx1_ASAP7_6t_fix 0 0 ;
  SIZE 0.864 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN L
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.268 0.516 0.576 0.588 ;
        RECT 0.504 0.108 0.576 0.588 ;
        RECT 0.356 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.288 0.516 0.36 0.588 ;
        RECT 0.396 0.108 0.468 0.18 ;
    END
  END L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 0.864 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 0.864 0.912 ;
        RECT 0.384 0.648 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 0.864 0.048 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.072 0.684 0.292 0.756 ;
      RECT 0.072 0.272 0.144 0.756 ;
      RECT 0.072 0.272 0.34 0.344 ;
  END
END TIELOx1_ASAP7_6t_fix

MACRO XNOR2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.228 0.252 2.136 0.324 ;
      LAYER M1 ;
        RECT 2.044 0.244 2.116 0.488 ;
        RECT 1.256 0.396 1.46 0.468 ;
        RECT 1.256 0.252 1.328 0.468 ;
        RECT 0.828 0.252 1.328 0.324 ;
        RECT 0.828 0.108 0.9 0.324 ;
        RECT 0.072 0.108 0.9 0.18 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V1 ;
        RECT 1.248 0.252 1.32 0.324 ;
        RECT 2.044 0.252 2.116 0.324 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 1.368 0.396 1.44 0.468 ;
        RECT 2.044 0.396 2.116 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 1.896 0.54 1.992 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.684 2.432 0.756 ;
        RECT 1.872 0.252 1.944 0.756 ;
        RECT 1.672 0.252 1.944 0.324 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.252 1.764 0.324 ;
        RECT 2.34 0.684 2.412 0.756 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.592 0.54 2.332 0.612 ;
      LAYER M1 ;
        RECT 2.232 0.54 2.38 0.612 ;
        RECT 2.232 0.384 2.304 0.612 ;
        RECT 0.612 0.396 0.944 0.468 ;
        RECT 0.612 0.396 0.684 0.62 ;
      LAYER V1 ;
        RECT 0.612 0.54 0.684 0.612 ;
        RECT 2.24 0.54 2.312 0.612 ;
      LAYER V0 ;
        RECT 0.852 0.396 0.924 0.468 ;
        RECT 2.232 0.404 2.304 0.476 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 0.772 0.684 0.92 0.756 ;
      RECT 0.848 0.54 0.92 0.756 ;
      RECT 0.848 0.54 1.656 0.612 ;
      RECT 1.584 0.396 1.656 0.612 ;
      RECT 1.584 0.396 1.764 0.468 ;
      RECT 0.376 0.684 0.54 0.756 ;
      RECT 0.468 0.252 0.54 0.756 ;
      RECT 0.468 0.252 0.704 0.324 ;
      RECT 2.284 0.108 2.432 0.18 ;
      RECT 1.784 0.108 1.98 0.18 ;
      RECT 1.024 0.108 1.548 0.18 ;
    LAYER M2 ;
      RECT 1.448 0.108 2.432 0.18 ;
      RECT 0.376 0.684 0.872 0.756 ;
    LAYER V1 ;
      RECT 2.34 0.108 2.412 0.18 ;
      RECT 1.836 0.108 1.908 0.18 ;
      RECT 1.468 0.108 1.54 0.18 ;
      RECT 0.78 0.684 0.852 0.756 ;
      RECT 0.396 0.684 0.468 0.756 ;
  END
END XNOR2x1_ASAP7_6t_fix

MACRO XNOR2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.552 0.54 1.78 0.612 ;
      LAYER M1 ;
        RECT 1.688 0.4 1.76 0.62 ;
        RECT 1.564 0.4 1.76 0.472 ;
        RECT 0.504 0.54 0.652 0.612 ;
        RECT 0.504 0.38 0.576 0.612 ;
      LAYER V1 ;
        RECT 0.572 0.54 0.644 0.612 ;
        RECT 1.688 0.54 1.76 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.4 0.576 0.472 ;
        RECT 1.584 0.4 1.656 0.472 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.684 1.516 0.756 ;
        RECT 1.368 0.396 1.44 0.756 ;
      LAYER V0 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 0.6 0.54 0.696 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 1.248 -0.048 1.344 0.216 ;
        RECT 0.384 -0.048 0.48 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.684 2.304 0.756 ;
        RECT 2.232 0.108 2.304 0.756 ;
        RECT 1.888 0.108 2.304 0.18 ;
      LAYER V0 ;
        RECT 1.908 0.684 1.98 0.756 ;
        RECT 1.908 0.108 1.98 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.908 0.252 1.98 0.488 ;
      RECT 1.692 0.252 1.98 0.324 ;
      RECT 1.188 0.108 1.26 0.612 ;
      RECT 0.288 0.108 0.36 0.584 ;
      RECT 0.288 0.108 1.568 0.18 ;
      RECT 0.072 0.684 0.252 0.756 ;
      RECT 0.072 0.232 0.144 0.756 ;
      RECT 0.712 0.252 0.92 0.324 ;
      RECT 0.396 0.684 0.92 0.756 ;
    LAYER M2 ;
      RECT 0.052 0.252 1.792 0.324 ;
    LAYER V1 ;
      RECT 1.7 0.252 1.772 0.324 ;
      RECT 0.828 0.252 0.9 0.324 ;
      RECT 0.072 0.252 0.144 0.324 ;
  END
END XNOR2x2_ASAP7_6t_fix

MACRO XNOR2xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.072 0.252 0.928 0.324 ;
      LAYER M1 ;
        RECT 1.292 0.396 1.512 0.468 ;
        RECT 1.44 0.252 1.512 0.468 ;
        RECT 0.828 0.252 1.512 0.324 ;
        RECT 0.072 0.684 0.22 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V1 ;
        RECT 0.072 0.252 0.144 0.324 ;
        RECT 0.836 0.252 0.908 0.324 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 1.368 0.396 1.44 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.54 0.576 0.612 ;
        RECT 0.504 0.108 0.576 0.612 ;
        RECT 0.428 0.108 0.576 0.18 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.464 0.54 1.56 0.912 ;
        RECT 0.6 0.648 0.696 0.912 ;
        RECT 0.168 0.648 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.248 -0.048 1.344 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.692 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.044 0.684 1.116 0.756 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.684 0.728 0.756 ;
      RECT 0.656 0.252 0.728 0.756 ;
      RECT 0.656 0.54 1.656 0.612 ;
      RECT 1.584 0.376 1.656 0.612 ;
      RECT 1.044 0.108 1.548 0.18 ;
  END
END XNOR2xp5_ASAP7_6t_fix

MACRO XOR2x1_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1_ASAP7_6t_fix 0 0 ;
  SIZE 2.592 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.88 0.54 2.108 0.612 ;
      LAYER M1 ;
        RECT 2.008 0.54 2.164 0.612 ;
        RECT 2.016 0.396 2.088 0.612 ;
        RECT 0.9 0.396 1.46 0.468 ;
        RECT 0.072 0.684 0.972 0.756 ;
        RECT 0.9 0.396 0.972 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V1 ;
        RECT 0.9 0.54 0.972 0.612 ;
        RECT 2.016 0.54 2.088 0.612 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 1.364 0.396 1.436 0.468 ;
        RECT 2.016 0.396 2.088 0.468 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.592 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.592 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
        RECT 2.34 0.828 2.412 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.592 0.048 ;
        RECT 1.896 -0.048 1.992 0.324 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
        RECT 0.168 -0.048 0.264 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
        RECT 2.34 -0.036 2.412 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.108 2.196 0.18 ;
        RECT 1.7 0.54 1.872 0.612 ;
        RECT 1.8 0.108 1.872 0.612 ;
      LAYER V0 ;
        RECT 1.044 0.108 1.116 0.18 ;
        RECT 1.692 0.108 1.764 0.18 ;
        RECT 1.72 0.54 1.792 0.612 ;
        RECT 2.124 0.108 2.196 0.18 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.452 0.252 2.304 0.324 ;
      LAYER M1 ;
        RECT 2.168 0.252 2.316 0.324 ;
        RECT 2.232 0.252 2.304 0.488 ;
        RECT 0.504 0.252 0.576 0.488 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V1 ;
        RECT 0.472 0.252 0.544 0.324 ;
        RECT 2.232 0.252 2.304 0.324 ;
      LAYER V0 ;
        RECT 0.504 0.396 0.576 0.468 ;
        RECT 2.232 0.396 2.304 0.468 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 1.044 0.684 2.432 0.756 ;
      RECT 1.044 0.592 1.116 0.756 ;
      RECT 0.664 0.54 0.828 0.612 ;
      RECT 0.756 0.108 0.828 0.612 ;
      RECT 1.56 0.252 1.632 0.48 ;
      RECT 0.756 0.252 1.632 0.324 ;
      RECT 0.368 0.108 0.828 0.18 ;
  END
END XOR2x1_ASAP7_6t_fix

MACRO XOR2x2_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x2_ASAP7_6t_fix 0 0 ;
  SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.308 0.396 1.48 0.468 ;
        RECT 1.408 0.108 1.48 0.468 ;
        RECT 1.288 0.108 1.48 0.18 ;
      LAYER V0 ;
        RECT 1.308 0.396 1.38 0.468 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.956 0.252 1.836 0.324 ;
      LAYER M1 ;
        RECT 1.584 0.396 1.836 0.468 ;
        RECT 1.764 0.108 1.836 0.468 ;
        RECT 1.644 0.108 1.836 0.18 ;
        RECT 0.616 0.252 1.036 0.324 ;
        RECT 0.488 0.396 0.688 0.468 ;
        RECT 0.616 0.252 0.688 0.468 ;
      LAYER V1 ;
        RECT 0.956 0.252 1.028 0.324 ;
        RECT 1.764 0.252 1.836 0.324 ;
      LAYER V0 ;
        RECT 0.508 0.396 0.58 0.468 ;
        RECT 1.612 0.396 1.684 0.468 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 2.376 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 2.376 0.912 ;
        RECT 2.112 0.54 2.208 0.912 ;
        RECT 1.68 0.54 1.776 0.912 ;
        RECT 1.248 0.648 1.344 0.912 ;
        RECT 0.384 0.54 0.48 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
        RECT 1.908 0.828 1.98 0.9 ;
        RECT 2.124 0.828 2.196 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 2.376 0.048 ;
        RECT 2.112 -0.048 2.208 0.324 ;
        RECT 1.68 -0.048 1.776 0.324 ;
        RECT 0.6 -0.048 0.696 0.324 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
        RECT 1.908 -0.036 1.98 0.036 ;
        RECT 2.124 -0.036 2.196 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.684 2.304 0.756 ;
        RECT 2.232 0.108 2.304 0.756 ;
        RECT 1.908 0.108 2.304 0.18 ;
        RECT 1.908 0.108 1.98 0.272 ;
      LAYER V0 ;
        RECT 1.908 0.684 1.98 0.756 ;
        RECT 1.908 0.18 1.98 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.308 0.54 1.98 0.612 ;
      RECT 1.908 0.388 1.98 0.612 ;
      RECT 1.908 0.388 2.112 0.46 ;
      RECT 0.316 0.684 1.568 0.756 ;
      RECT 1.136 0.232 1.208 0.756 ;
      RECT 0.316 0.376 0.388 0.756 ;
      RECT 0.796 0.54 0.944 0.612 ;
      RECT 0.396 0.108 0.92 0.18 ;
      RECT 0.072 0.54 0.216 0.612 ;
    LAYER M2 ;
      RECT 0.136 0.54 1.388 0.612 ;
    LAYER V1 ;
      RECT 1.316 0.54 1.388 0.612 ;
      RECT 0.828 0.54 0.9 0.612 ;
      RECT 0.136 0.54 0.208 0.612 ;
  END
END XOR2x2_ASAP7_6t_fix

MACRO XOR2xp5_ASAP7_6t_fix
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2xp5_ASAP7_6t_fix 0 0 ;
  SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.412 1.44 0.484 ;
        RECT 0.844 0.536 1.172 0.608 ;
        RECT 1.1 0.412 1.172 0.608 ;
        RECT 0.072 0.684 0.916 0.756 ;
        RECT 0.844 0.536 0.916 0.756 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.756 ;
      LAYER V0 ;
        RECT 0.072 0.396 0.144 0.468 ;
        RECT 1.368 0.412 1.44 0.484 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.332 0.576 0.404 ;
        RECT 0.288 0.252 0.504 0.612 ;
      LAYER V0 ;
        RECT 0.504 0.332 0.576 0.404 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.828 1.944 0.9 ;
      LAYER LISD ;
        RECT 0 0.816 1.944 0.912 ;
        RECT 1.248 0.54 1.344 0.912 ;
        RECT 0.168 0.54 0.264 0.912 ;
      LAYER V0 ;
        RECT 0.18 0.828 0.252 0.9 ;
        RECT 0.396 0.828 0.468 0.9 ;
        RECT 0.612 0.828 0.684 0.9 ;
        RECT 0.828 0.828 0.9 0.9 ;
        RECT 1.044 0.828 1.116 0.9 ;
        RECT 1.26 0.828 1.332 0.9 ;
        RECT 1.476 0.828 1.548 0.9 ;
        RECT 1.692 0.828 1.764 0.9 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
      LAYER LISD ;
        RECT 0 -0.048 1.944 0.048 ;
        RECT 1.464 -0.048 1.56 0.324 ;
        RECT 0.6 -0.048 0.696 0.216 ;
        RECT 0.168 -0.048 0.264 0.216 ;
      LAYER V0 ;
        RECT 0.18 -0.036 0.252 0.036 ;
        RECT 0.396 -0.036 0.468 0.036 ;
        RECT 0.612 -0.036 0.684 0.036 ;
        RECT 0.828 -0.036 0.9 0.036 ;
        RECT 1.044 -0.036 1.116 0.036 ;
        RECT 1.26 -0.036 1.332 0.036 ;
        RECT 1.476 -0.036 1.548 0.036 ;
        RECT 1.692 -0.036 1.764 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.684 1.872 0.756 ;
        RECT 1.8 0.108 1.872 0.756 ;
        RECT 1.26 0.108 1.872 0.18 ;
      LAYER V0 ;
        RECT 1.26 0.108 1.332 0.18 ;
        RECT 1.692 0.684 1.764 0.756 ;
        RECT 1.692 0.108 1.764 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.608 0.54 0.756 0.612 ;
      RECT 0.684 0.108 0.756 0.612 ;
      RECT 1.584 0.252 1.656 0.488 ;
      RECT 0.684 0.252 1.656 0.324 ;
      RECT 0.396 0.108 0.756 0.18 ;
      RECT 1.044 0.684 1.548 0.756 ;
  END
END XOR2xp5_ASAP7_6t_fix

END LIBRARY
